// Benchmark "cir1_cir2_miter" written by ABC on Thu Jul 13 12:02:42 2023

module cir1_cir2_miter ( 
    controlPi_0_0, controlPi_0_1, controlPi_0_2, controlPi_0_3,
    controlPi_0_4, controlPi_0_5, controlPi_0_6, controlPi_0_7,
    controlPi_1_0, controlPi_1_1, controlPi_1_2, controlPi_1_3,
    controlPi_1_4, controlPi_1_5, controlPi_1_6, controlPi_1_7,
    controlPi_2_0, controlPi_2_1, controlPi_2_2, controlPi_2_3,
    controlPi_2_4, controlPi_2_5, controlPi_2_6, controlPi_2_7,
    controlPi_3_0, controlPi_3_1, controlPi_3_2, controlPi_3_3,
    controlPi_3_4, controlPi_3_5, controlPi_3_6, controlPi_3_7,
    controlPi_4_0, controlPi_4_1, controlPi_4_2, controlPi_4_3,
    controlPi_4_4, controlPi_4_5, controlPi_4_6, controlPi_4_7,
    controlPi_5_0, controlPi_5_1, controlPi_5_2, controlPi_5_3,
    controlPi_5_4, controlPi_5_5, controlPi_5_6, controlPi_5_7,
    controlPi_6_0, controlPi_6_1, controlPi_6_2, controlPi_6_3,
    controlPi_6_4, controlPi_6_5, controlPi_6_6, controlPi_6_7,
    controlPi_7_0, controlPi_7_1, controlPi_7_2, controlPi_7_3,
    controlPi_7_4, controlPi_7_5, controlPi_7_6, controlPi_7_7,
    controlPi_8_0, controlPi_8_1, controlPi_8_2, controlPi_8_3,
    controlPi_8_4, controlPi_8_5, controlPi_8_6, controlPi_8_7,
    controlPi_9_0, controlPi_9_1, controlPi_9_2, controlPi_9_3,
    controlPi_9_4, controlPi_9_5, controlPi_9_6, controlPi_9_7,
    controlPi_10_0, controlPi_10_1, controlPi_10_2, controlPi_10_3,
    controlPi_10_4, controlPi_10_5, controlPi_10_6, controlPi_10_7,
    controlPi_11_0, controlPi_11_1, controlPi_11_2, controlPi_11_3,
    controlPi_11_4, controlPi_11_5, controlPi_11_6, controlPi_11_7,
    controlPi_12_0, controlPi_12_1, controlPi_12_2, controlPi_12_3,
    controlPi_12_4, controlPi_12_5, controlPi_12_6, controlPi_12_7,
    controlPi_13_0, controlPi_13_1, controlPi_13_2, controlPi_13_3,
    controlPi_13_4, controlPi_13_5, controlPi_13_6, controlPi_13_7,
    controlPi_14_0, controlPi_14_1, controlPi_14_2, controlPi_14_3,
    controlPi_14_4, controlPi_14_5, controlPi_14_6, controlPi_14_7,
    controlPi_15_0, controlPi_15_1, controlPi_15_2, controlPi_15_3,
    controlPi_15_4, controlPi_15_5, controlPi_15_6, controlPi_15_7,
    controlPi_16_0, controlPi_16_1, controlPi_16_2, controlPi_16_3,
    controlPi_16_4, controlPi_16_5, controlPi_16_6, controlPi_16_7,
    controlPi_17_0, controlPi_17_1, controlPi_17_2, controlPi_17_3,
    controlPi_17_4, controlPi_17_5, controlPi_17_6, controlPi_17_7,
    controlPi_18_0, controlPi_18_1, controlPi_18_2, controlPi_18_3,
    controlPi_18_4, controlPi_18_5, controlPi_18_6, controlPi_18_7,
    controlPi_19_0, controlPi_19_1, controlPi_19_2, controlPi_19_3,
    controlPi_19_4, controlPi_19_5, controlPi_19_6, controlPi_19_7,
    controlPi_20_0, controlPi_20_1, controlPi_20_2, controlPi_20_3,
    controlPi_20_4, controlPi_20_5, controlPi_20_6, controlPi_20_7,
    controlPi_21_0, controlPi_21_1, controlPi_21_2, controlPi_21_3,
    controlPi_21_4, controlPi_21_5, controlPi_21_6, controlPi_21_7,
    controlPi_22_0, controlPi_22_1, controlPi_22_2, controlPi_22_3,
    controlPi_22_4, controlPi_22_5, controlPi_22_6, controlPi_22_7,
    controlPi_23_0, controlPi_23_1, controlPi_23_2, controlPi_23_3,
    controlPi_23_4, controlPi_23_5, controlPi_23_6, controlPi_23_7,
    controlPi_24_0, controlPi_24_1, controlPi_24_2, controlPi_24_3,
    controlPi_24_4, controlPi_24_5, controlPi_24_6, controlPi_24_7,
    controlPi_25_0, controlPi_25_1, controlPi_25_2, controlPi_25_3,
    controlPi_25_4, controlPi_25_5, controlPi_25_6, controlPi_25_7,
    controlPi_26_0, controlPi_26_1, controlPi_26_2, controlPi_26_3,
    controlPi_26_4, controlPi_26_5, controlPi_26_6, controlPi_26_7,
    controlPi_27_0, controlPi_27_1, controlPi_27_2, controlPi_27_3,
    controlPi_27_4, controlPi_27_5, controlPi_27_6, controlPi_27_7,
    controlPi_28_0, controlPi_28_1, controlPi_28_2, controlPi_28_3,
    controlPi_28_4, controlPi_28_5, controlPi_28_6, controlPi_28_7,
    controlPi_29_0, controlPi_29_1, controlPi_29_2, controlPi_29_3,
    controlPi_29_4, controlPi_29_5, controlPi_29_6, controlPi_29_7,
    controlPi_30_0, controlPi_30_1, controlPi_30_2, controlPi_30_3,
    controlPi_30_4, controlPi_30_5, controlPi_30_6, controlPi_30_7,
    controlPi_31_0, controlPi_31_1, controlPi_31_2, controlPi_31_3,
    controlPi_31_4, controlPi_31_5, controlPi_31_6, controlPi_31_7,
    controlPi_32_0, controlPi_32_1, controlPi_32_2, controlPi_32_3,
    controlPi_32_4, controlPi_32_5, controlPi_32_6, controlPi_32_7,
    controlPi_33_0, controlPi_33_1, controlPi_33_2, controlPi_33_3,
    controlPi_33_4, controlPi_33_5, controlPi_33_6, controlPi_33_7,
    controlPi_34_0, controlPi_34_1, controlPi_34_2, controlPi_34_3,
    controlPi_34_4, controlPi_34_5, controlPi_34_6, controlPi_34_7,
    controlPi_35_0, controlPi_35_1, controlPi_35_2, controlPi_35_3,
    controlPi_35_4, controlPi_35_5, controlPi_35_6, controlPi_35_7,
    controlPi_36_0, controlPi_36_1, controlPi_36_2, controlPi_36_3,
    controlPi_36_4, controlPi_36_5, controlPi_36_6, controlPi_36_7,
    controlPi_37_0, controlPi_37_1, controlPi_37_2, controlPi_37_3,
    controlPi_37_4, controlPi_37_5, controlPi_37_6, controlPi_37_7,
    controlPi_38_0, controlPi_38_1, controlPi_38_2, controlPi_38_3,
    controlPi_38_4, controlPi_38_5, controlPi_38_6, controlPi_38_7,
    controlPi_39_0, controlPi_39_1, controlPi_39_2, controlPi_39_3,
    controlPi_39_4, controlPi_39_5, controlPi_39_6, controlPi_39_7,
    controlPi_40_0, controlPi_40_1, controlPi_40_2, controlPi_40_3,
    controlPi_40_4, controlPi_40_5, controlPi_40_6, controlPi_40_7,
    controlPi_41_0, controlPi_41_1, controlPi_41_2, controlPi_41_3,
    controlPi_41_4, controlPi_41_5, controlPi_41_6, controlPi_41_7,
    controlPi_42_0, controlPi_42_1, controlPi_42_2, controlPi_42_3,
    controlPi_42_4, controlPi_42_5, controlPi_42_6, controlPi_42_7,
    controlPi_43_0, controlPi_43_1, controlPi_43_2, controlPi_43_3,
    controlPi_43_4, controlPi_43_5, controlPi_43_6, controlPi_43_7,
    controlPi_44_0, controlPi_44_1, controlPi_44_2, controlPi_44_3,
    controlPi_44_4, controlPi_44_5, controlPi_44_6, controlPi_44_7,
    controlPi_45_0, controlPi_45_1, controlPi_45_2, controlPi_45_3,
    controlPi_45_4, controlPi_45_5, controlPi_45_6, controlPi_45_7,
    controlPi_46_0, controlPi_46_1, controlPi_46_2, controlPi_46_3,
    controlPi_46_4, controlPi_46_5, controlPi_46_6, controlPi_46_7,
    controlPi_47_0, controlPi_47_1, controlPi_47_2, controlPi_47_3,
    controlPi_47_4, controlPi_47_5, controlPi_47_6, controlPi_47_7,
    controlPi_48_0, controlPi_48_1, controlPi_48_2, controlPi_48_3,
    controlPi_48_4, controlPi_48_5, controlPi_48_6, controlPi_48_7,
    controlPi_49_0, controlPi_49_1, controlPi_49_2, controlPi_49_3,
    controlPi_49_4, controlPi_49_5, controlPi_49_6, controlPi_49_7,
    controlPi_50_0, controlPi_50_1, controlPi_50_2, controlPi_50_3,
    controlPi_50_4, controlPi_50_5, controlPi_50_6, controlPi_50_7,
    controlPi_51_0, controlPi_51_1, controlPi_51_2, controlPi_51_3,
    controlPi_51_4, controlPi_51_5, controlPi_51_6, controlPi_51_7,
    controlPi_52_0, controlPi_52_1, controlPi_52_2, controlPi_52_3,
    controlPi_52_4, controlPi_52_5, controlPi_52_6, controlPi_52_7,
    controlPi_53_0, controlPi_53_1, controlPi_53_2, controlPi_53_3,
    controlPi_53_4, controlPi_53_5, controlPi_53_6, controlPi_53_7,
    controlPi_54_0, controlPi_54_1, controlPi_54_2, controlPi_54_3,
    controlPi_54_4, controlPi_54_5, controlPi_54_6, controlPi_54_7,
    controlPi_55_0, controlPi_55_1, controlPi_55_2, controlPi_55_3,
    controlPi_55_4, controlPi_55_5, controlPi_55_6, controlPi_55_7,
    controlPi_56_0, controlPi_56_1, controlPi_56_2, controlPi_56_3,
    controlPi_56_4, controlPi_56_5, controlPi_56_6, controlPi_56_7,
    controlPi_57_0, controlPi_57_1, controlPi_57_2, controlPi_57_3,
    controlPi_57_4, controlPi_57_5, controlPi_57_6, controlPi_57_7,
    controlPi_58_0, controlPi_58_1, controlPi_58_2, controlPi_58_3,
    controlPi_58_4, controlPi_58_5, controlPi_58_6, controlPi_58_7,
    controlPi_59_0, controlPi_59_1, controlPi_59_2, controlPi_59_3,
    controlPi_59_4, controlPi_59_5, controlPi_59_6, controlPi_59_7,
    controlPi_60_0, controlPi_60_1, controlPi_60_2, controlPi_60_3,
    controlPi_60_4, controlPi_60_5, controlPi_60_6, controlPi_60_7,
    controlPi_61_0, controlPi_61_1, controlPi_61_2, controlPi_61_3,
    controlPi_61_4, controlPi_61_5, controlPi_61_6, controlPi_61_7,
    controlPi_62_0, controlPi_62_1, controlPi_62_2, controlPi_62_3,
    controlPi_62_4, controlPi_62_5, controlPi_62_6, controlPi_62_7,
    controlPi_63_0, controlPi_63_1, controlPi_63_2, controlPi_63_3,
    controlPi_63_4, controlPi_63_5, controlPi_63_6, controlPi_63_7,
    controlPi_64_0, controlPi_64_1, controlPi_64_2, controlPi_64_3,
    controlPi_64_4, controlPi_64_5, controlPi_64_6, controlPi_64_7,
    controlPi_65_0, controlPi_65_1, controlPi_65_2, controlPi_65_3,
    controlPi_65_4, controlPi_65_5, controlPi_65_6, controlPi_65_7,
    controlPi_66_0, controlPi_66_1, controlPi_66_2, controlPi_66_3,
    controlPi_66_4, controlPi_66_5, controlPi_66_6, controlPi_66_7,
    controlPi_67_0, controlPi_67_1, controlPi_67_2, controlPi_67_3,
    controlPi_67_4, controlPi_67_5, controlPi_67_6, controlPi_67_7,
    controlPi_68_0, controlPi_68_1, controlPi_68_2, controlPi_68_3,
    controlPi_68_4, controlPi_68_5, controlPi_68_6, controlPi_68_7,
    controlPi_69_0, controlPi_69_1, controlPi_69_2, controlPi_69_3,
    controlPi_69_4, controlPi_69_5, controlPi_69_6, controlPi_69_7,
    controlPi_70_0, controlPi_70_1, controlPi_70_2, controlPi_70_3,
    controlPi_70_4, controlPi_70_5, controlPi_70_6, controlPi_70_7,
    controlPi_71_0, controlPi_71_1, controlPi_71_2, controlPi_71_3,
    controlPi_71_4, controlPi_71_5, controlPi_71_6, controlPi_71_7,
    controlPi_72_0, controlPi_72_1, controlPi_72_2, controlPi_72_3,
    controlPi_72_4, controlPi_72_5, controlPi_72_6, controlPi_72_7,
    controlPi_73_0, controlPi_73_1, controlPi_73_2, controlPi_73_3,
    controlPi_73_4, controlPi_73_5, controlPi_73_6, controlPi_73_7,
    controlPi_74_0, controlPi_74_1, controlPi_74_2, controlPi_74_3,
    controlPi_74_4, controlPi_74_5, controlPi_74_6, controlPi_74_7,
    controlPi_75_0, controlPi_75_1, controlPi_75_2, controlPi_75_3,
    controlPi_75_4, controlPi_75_5, controlPi_75_6, controlPi_75_7,
    controlPi_76_0, controlPi_76_1, controlPi_76_2, controlPi_76_3,
    controlPi_76_4, controlPi_76_5, controlPi_76_6, controlPi_76_7,
    controlPi_77_0, controlPi_77_1, controlPi_77_2, controlPi_77_3,
    controlPi_77_4, controlPi_77_5, controlPi_77_6, controlPi_77_7,
    controlPi_78_0, controlPi_78_1, controlPi_78_2, controlPi_78_3,
    controlPi_78_4, controlPi_78_5, controlPi_78_6, controlPi_78_7,
    controlPi_79_0, controlPi_79_1, controlPi_79_2, controlPi_79_3,
    controlPi_79_4, controlPi_79_5, controlPi_79_6, controlPi_79_7,
    controlPi_80_0, controlPi_80_1, controlPi_80_2, controlPi_80_3,
    controlPi_80_4, controlPi_80_5, controlPi_80_6, controlPi_80_7,
    controlPi_81_0, controlPi_81_1, controlPi_81_2, controlPi_81_3,
    controlPi_81_4, controlPi_81_5, controlPi_81_6, controlPi_81_7,
    controlPi_82_0, controlPi_82_1, controlPi_82_2, controlPi_82_3,
    controlPi_82_4, controlPi_82_5, controlPi_82_6, controlPi_82_7,
    controlPi_83_0, controlPi_83_1, controlPi_83_2, controlPi_83_3,
    controlPi_83_4, controlPi_83_5, controlPi_83_6, controlPi_83_7,
    controlPi_84_0, controlPi_84_1, controlPi_84_2, controlPi_84_3,
    controlPi_84_4, controlPi_84_5, controlPi_84_6, controlPi_84_7,
    controlPi_85_0, controlPi_85_1, controlPi_85_2, controlPi_85_3,
    controlPi_85_4, controlPi_85_5, controlPi_85_6, controlPi_85_7,
    n2_ntk1, n11_ntk1, n13_ntk1, n16_ntk1, n21_ntk1, n45_ntk1, n46_ntk1,
    n55_ntk1, n74_ntk1, n75_ntk1, n81_ntk1, n84_ntk1, n85_ntk1, n93_ntk1,
    n96_ntk1, n98_ntk1, n101_ntk1, n111_ntk1, n128_ntk1, n131_ntk1,
    n134_ntk1, n139_ntk1, n153_ntk1, n159_ntk1, n177_ntk1, n199_ntk1,
    n206_ntk1, n211_ntk1, n216_ntk1, n223_ntk1, n243_ntk1, n264_ntk1,
    n266_ntk1, n280_ntk1, n282_ntk1, n287_ntk1, n290_ntk1, n309_ntk1,
    n336_ntk1, n346_ntk1, n349_ntk1, n360_ntk1, n368_ntk1, n369_ntk1,
    n377_ntk1, n388_ntk1, n394_ntk1, n409_ntk1, n428_ntk1, n435_ntk1,
    n447_ntk1, n454_ntk1, n457_ntk1, n468_ntk1, n471_ntk1, n481_ntk1,
    n494_ntk1, n500_ntk1, n507_ntk1, n511_ntk1, n519_ntk1, n525_ntk1,
    n557_ntk1, n561_ntk1, n569_ntk1, n571_ntk1, n575_ntk1, n581_ntk1,
    n582_ntk1, n583_ntk1, n587_ntk1, n600_ntk1, n603_ntk1, n609_ntk1,
    n613_ntk1, n614_ntk1, n616_ntk1, n646_ntk1, n659_ntk1, n661_ntk1,
    n664_ntk1, n673_ntk1,
    miter  );
  input  controlPi_0_0, controlPi_0_1, controlPi_0_2, controlPi_0_3,
    controlPi_0_4, controlPi_0_5, controlPi_0_6, controlPi_0_7,
    controlPi_1_0, controlPi_1_1, controlPi_1_2, controlPi_1_3,
    controlPi_1_4, controlPi_1_5, controlPi_1_6, controlPi_1_7,
    controlPi_2_0, controlPi_2_1, controlPi_2_2, controlPi_2_3,
    controlPi_2_4, controlPi_2_5, controlPi_2_6, controlPi_2_7,
    controlPi_3_0, controlPi_3_1, controlPi_3_2, controlPi_3_3,
    controlPi_3_4, controlPi_3_5, controlPi_3_6, controlPi_3_7,
    controlPi_4_0, controlPi_4_1, controlPi_4_2, controlPi_4_3,
    controlPi_4_4, controlPi_4_5, controlPi_4_6, controlPi_4_7,
    controlPi_5_0, controlPi_5_1, controlPi_5_2, controlPi_5_3,
    controlPi_5_4, controlPi_5_5, controlPi_5_6, controlPi_5_7,
    controlPi_6_0, controlPi_6_1, controlPi_6_2, controlPi_6_3,
    controlPi_6_4, controlPi_6_5, controlPi_6_6, controlPi_6_7,
    controlPi_7_0, controlPi_7_1, controlPi_7_2, controlPi_7_3,
    controlPi_7_4, controlPi_7_5, controlPi_7_6, controlPi_7_7,
    controlPi_8_0, controlPi_8_1, controlPi_8_2, controlPi_8_3,
    controlPi_8_4, controlPi_8_5, controlPi_8_6, controlPi_8_7,
    controlPi_9_0, controlPi_9_1, controlPi_9_2, controlPi_9_3,
    controlPi_9_4, controlPi_9_5, controlPi_9_6, controlPi_9_7,
    controlPi_10_0, controlPi_10_1, controlPi_10_2, controlPi_10_3,
    controlPi_10_4, controlPi_10_5, controlPi_10_6, controlPi_10_7,
    controlPi_11_0, controlPi_11_1, controlPi_11_2, controlPi_11_3,
    controlPi_11_4, controlPi_11_5, controlPi_11_6, controlPi_11_7,
    controlPi_12_0, controlPi_12_1, controlPi_12_2, controlPi_12_3,
    controlPi_12_4, controlPi_12_5, controlPi_12_6, controlPi_12_7,
    controlPi_13_0, controlPi_13_1, controlPi_13_2, controlPi_13_3,
    controlPi_13_4, controlPi_13_5, controlPi_13_6, controlPi_13_7,
    controlPi_14_0, controlPi_14_1, controlPi_14_2, controlPi_14_3,
    controlPi_14_4, controlPi_14_5, controlPi_14_6, controlPi_14_7,
    controlPi_15_0, controlPi_15_1, controlPi_15_2, controlPi_15_3,
    controlPi_15_4, controlPi_15_5, controlPi_15_6, controlPi_15_7,
    controlPi_16_0, controlPi_16_1, controlPi_16_2, controlPi_16_3,
    controlPi_16_4, controlPi_16_5, controlPi_16_6, controlPi_16_7,
    controlPi_17_0, controlPi_17_1, controlPi_17_2, controlPi_17_3,
    controlPi_17_4, controlPi_17_5, controlPi_17_6, controlPi_17_7,
    controlPi_18_0, controlPi_18_1, controlPi_18_2, controlPi_18_3,
    controlPi_18_4, controlPi_18_5, controlPi_18_6, controlPi_18_7,
    controlPi_19_0, controlPi_19_1, controlPi_19_2, controlPi_19_3,
    controlPi_19_4, controlPi_19_5, controlPi_19_6, controlPi_19_7,
    controlPi_20_0, controlPi_20_1, controlPi_20_2, controlPi_20_3,
    controlPi_20_4, controlPi_20_5, controlPi_20_6, controlPi_20_7,
    controlPi_21_0, controlPi_21_1, controlPi_21_2, controlPi_21_3,
    controlPi_21_4, controlPi_21_5, controlPi_21_6, controlPi_21_7,
    controlPi_22_0, controlPi_22_1, controlPi_22_2, controlPi_22_3,
    controlPi_22_4, controlPi_22_5, controlPi_22_6, controlPi_22_7,
    controlPi_23_0, controlPi_23_1, controlPi_23_2, controlPi_23_3,
    controlPi_23_4, controlPi_23_5, controlPi_23_6, controlPi_23_7,
    controlPi_24_0, controlPi_24_1, controlPi_24_2, controlPi_24_3,
    controlPi_24_4, controlPi_24_5, controlPi_24_6, controlPi_24_7,
    controlPi_25_0, controlPi_25_1, controlPi_25_2, controlPi_25_3,
    controlPi_25_4, controlPi_25_5, controlPi_25_6, controlPi_25_7,
    controlPi_26_0, controlPi_26_1, controlPi_26_2, controlPi_26_3,
    controlPi_26_4, controlPi_26_5, controlPi_26_6, controlPi_26_7,
    controlPi_27_0, controlPi_27_1, controlPi_27_2, controlPi_27_3,
    controlPi_27_4, controlPi_27_5, controlPi_27_6, controlPi_27_7,
    controlPi_28_0, controlPi_28_1, controlPi_28_2, controlPi_28_3,
    controlPi_28_4, controlPi_28_5, controlPi_28_6, controlPi_28_7,
    controlPi_29_0, controlPi_29_1, controlPi_29_2, controlPi_29_3,
    controlPi_29_4, controlPi_29_5, controlPi_29_6, controlPi_29_7,
    controlPi_30_0, controlPi_30_1, controlPi_30_2, controlPi_30_3,
    controlPi_30_4, controlPi_30_5, controlPi_30_6, controlPi_30_7,
    controlPi_31_0, controlPi_31_1, controlPi_31_2, controlPi_31_3,
    controlPi_31_4, controlPi_31_5, controlPi_31_6, controlPi_31_7,
    controlPi_32_0, controlPi_32_1, controlPi_32_2, controlPi_32_3,
    controlPi_32_4, controlPi_32_5, controlPi_32_6, controlPi_32_7,
    controlPi_33_0, controlPi_33_1, controlPi_33_2, controlPi_33_3,
    controlPi_33_4, controlPi_33_5, controlPi_33_6, controlPi_33_7,
    controlPi_34_0, controlPi_34_1, controlPi_34_2, controlPi_34_3,
    controlPi_34_4, controlPi_34_5, controlPi_34_6, controlPi_34_7,
    controlPi_35_0, controlPi_35_1, controlPi_35_2, controlPi_35_3,
    controlPi_35_4, controlPi_35_5, controlPi_35_6, controlPi_35_7,
    controlPi_36_0, controlPi_36_1, controlPi_36_2, controlPi_36_3,
    controlPi_36_4, controlPi_36_5, controlPi_36_6, controlPi_36_7,
    controlPi_37_0, controlPi_37_1, controlPi_37_2, controlPi_37_3,
    controlPi_37_4, controlPi_37_5, controlPi_37_6, controlPi_37_7,
    controlPi_38_0, controlPi_38_1, controlPi_38_2, controlPi_38_3,
    controlPi_38_4, controlPi_38_5, controlPi_38_6, controlPi_38_7,
    controlPi_39_0, controlPi_39_1, controlPi_39_2, controlPi_39_3,
    controlPi_39_4, controlPi_39_5, controlPi_39_6, controlPi_39_7,
    controlPi_40_0, controlPi_40_1, controlPi_40_2, controlPi_40_3,
    controlPi_40_4, controlPi_40_5, controlPi_40_6, controlPi_40_7,
    controlPi_41_0, controlPi_41_1, controlPi_41_2, controlPi_41_3,
    controlPi_41_4, controlPi_41_5, controlPi_41_6, controlPi_41_7,
    controlPi_42_0, controlPi_42_1, controlPi_42_2, controlPi_42_3,
    controlPi_42_4, controlPi_42_5, controlPi_42_6, controlPi_42_7,
    controlPi_43_0, controlPi_43_1, controlPi_43_2, controlPi_43_3,
    controlPi_43_4, controlPi_43_5, controlPi_43_6, controlPi_43_7,
    controlPi_44_0, controlPi_44_1, controlPi_44_2, controlPi_44_3,
    controlPi_44_4, controlPi_44_5, controlPi_44_6, controlPi_44_7,
    controlPi_45_0, controlPi_45_1, controlPi_45_2, controlPi_45_3,
    controlPi_45_4, controlPi_45_5, controlPi_45_6, controlPi_45_7,
    controlPi_46_0, controlPi_46_1, controlPi_46_2, controlPi_46_3,
    controlPi_46_4, controlPi_46_5, controlPi_46_6, controlPi_46_7,
    controlPi_47_0, controlPi_47_1, controlPi_47_2, controlPi_47_3,
    controlPi_47_4, controlPi_47_5, controlPi_47_6, controlPi_47_7,
    controlPi_48_0, controlPi_48_1, controlPi_48_2, controlPi_48_3,
    controlPi_48_4, controlPi_48_5, controlPi_48_6, controlPi_48_7,
    controlPi_49_0, controlPi_49_1, controlPi_49_2, controlPi_49_3,
    controlPi_49_4, controlPi_49_5, controlPi_49_6, controlPi_49_7,
    controlPi_50_0, controlPi_50_1, controlPi_50_2, controlPi_50_3,
    controlPi_50_4, controlPi_50_5, controlPi_50_6, controlPi_50_7,
    controlPi_51_0, controlPi_51_1, controlPi_51_2, controlPi_51_3,
    controlPi_51_4, controlPi_51_5, controlPi_51_6, controlPi_51_7,
    controlPi_52_0, controlPi_52_1, controlPi_52_2, controlPi_52_3,
    controlPi_52_4, controlPi_52_5, controlPi_52_6, controlPi_52_7,
    controlPi_53_0, controlPi_53_1, controlPi_53_2, controlPi_53_3,
    controlPi_53_4, controlPi_53_5, controlPi_53_6, controlPi_53_7,
    controlPi_54_0, controlPi_54_1, controlPi_54_2, controlPi_54_3,
    controlPi_54_4, controlPi_54_5, controlPi_54_6, controlPi_54_7,
    controlPi_55_0, controlPi_55_1, controlPi_55_2, controlPi_55_3,
    controlPi_55_4, controlPi_55_5, controlPi_55_6, controlPi_55_7,
    controlPi_56_0, controlPi_56_1, controlPi_56_2, controlPi_56_3,
    controlPi_56_4, controlPi_56_5, controlPi_56_6, controlPi_56_7,
    controlPi_57_0, controlPi_57_1, controlPi_57_2, controlPi_57_3,
    controlPi_57_4, controlPi_57_5, controlPi_57_6, controlPi_57_7,
    controlPi_58_0, controlPi_58_1, controlPi_58_2, controlPi_58_3,
    controlPi_58_4, controlPi_58_5, controlPi_58_6, controlPi_58_7,
    controlPi_59_0, controlPi_59_1, controlPi_59_2, controlPi_59_3,
    controlPi_59_4, controlPi_59_5, controlPi_59_6, controlPi_59_7,
    controlPi_60_0, controlPi_60_1, controlPi_60_2, controlPi_60_3,
    controlPi_60_4, controlPi_60_5, controlPi_60_6, controlPi_60_7,
    controlPi_61_0, controlPi_61_1, controlPi_61_2, controlPi_61_3,
    controlPi_61_4, controlPi_61_5, controlPi_61_6, controlPi_61_7,
    controlPi_62_0, controlPi_62_1, controlPi_62_2, controlPi_62_3,
    controlPi_62_4, controlPi_62_5, controlPi_62_6, controlPi_62_7,
    controlPi_63_0, controlPi_63_1, controlPi_63_2, controlPi_63_3,
    controlPi_63_4, controlPi_63_5, controlPi_63_6, controlPi_63_7,
    controlPi_64_0, controlPi_64_1, controlPi_64_2, controlPi_64_3,
    controlPi_64_4, controlPi_64_5, controlPi_64_6, controlPi_64_7,
    controlPi_65_0, controlPi_65_1, controlPi_65_2, controlPi_65_3,
    controlPi_65_4, controlPi_65_5, controlPi_65_6, controlPi_65_7,
    controlPi_66_0, controlPi_66_1, controlPi_66_2, controlPi_66_3,
    controlPi_66_4, controlPi_66_5, controlPi_66_6, controlPi_66_7,
    controlPi_67_0, controlPi_67_1, controlPi_67_2, controlPi_67_3,
    controlPi_67_4, controlPi_67_5, controlPi_67_6, controlPi_67_7,
    controlPi_68_0, controlPi_68_1, controlPi_68_2, controlPi_68_3,
    controlPi_68_4, controlPi_68_5, controlPi_68_6, controlPi_68_7,
    controlPi_69_0, controlPi_69_1, controlPi_69_2, controlPi_69_3,
    controlPi_69_4, controlPi_69_5, controlPi_69_6, controlPi_69_7,
    controlPi_70_0, controlPi_70_1, controlPi_70_2, controlPi_70_3,
    controlPi_70_4, controlPi_70_5, controlPi_70_6, controlPi_70_7,
    controlPi_71_0, controlPi_71_1, controlPi_71_2, controlPi_71_3,
    controlPi_71_4, controlPi_71_5, controlPi_71_6, controlPi_71_7,
    controlPi_72_0, controlPi_72_1, controlPi_72_2, controlPi_72_3,
    controlPi_72_4, controlPi_72_5, controlPi_72_6, controlPi_72_7,
    controlPi_73_0, controlPi_73_1, controlPi_73_2, controlPi_73_3,
    controlPi_73_4, controlPi_73_5, controlPi_73_6, controlPi_73_7,
    controlPi_74_0, controlPi_74_1, controlPi_74_2, controlPi_74_3,
    controlPi_74_4, controlPi_74_5, controlPi_74_6, controlPi_74_7,
    controlPi_75_0, controlPi_75_1, controlPi_75_2, controlPi_75_3,
    controlPi_75_4, controlPi_75_5, controlPi_75_6, controlPi_75_7,
    controlPi_76_0, controlPi_76_1, controlPi_76_2, controlPi_76_3,
    controlPi_76_4, controlPi_76_5, controlPi_76_6, controlPi_76_7,
    controlPi_77_0, controlPi_77_1, controlPi_77_2, controlPi_77_3,
    controlPi_77_4, controlPi_77_5, controlPi_77_6, controlPi_77_7,
    controlPi_78_0, controlPi_78_1, controlPi_78_2, controlPi_78_3,
    controlPi_78_4, controlPi_78_5, controlPi_78_6, controlPi_78_7,
    controlPi_79_0, controlPi_79_1, controlPi_79_2, controlPi_79_3,
    controlPi_79_4, controlPi_79_5, controlPi_79_6, controlPi_79_7,
    controlPi_80_0, controlPi_80_1, controlPi_80_2, controlPi_80_3,
    controlPi_80_4, controlPi_80_5, controlPi_80_6, controlPi_80_7,
    controlPi_81_0, controlPi_81_1, controlPi_81_2, controlPi_81_3,
    controlPi_81_4, controlPi_81_5, controlPi_81_6, controlPi_81_7,
    controlPi_82_0, controlPi_82_1, controlPi_82_2, controlPi_82_3,
    controlPi_82_4, controlPi_82_5, controlPi_82_6, controlPi_82_7,
    controlPi_83_0, controlPi_83_1, controlPi_83_2, controlPi_83_3,
    controlPi_83_4, controlPi_83_5, controlPi_83_6, controlPi_83_7,
    controlPi_84_0, controlPi_84_1, controlPi_84_2, controlPi_84_3,
    controlPi_84_4, controlPi_84_5, controlPi_84_6, controlPi_84_7,
    controlPi_85_0, controlPi_85_1, controlPi_85_2, controlPi_85_3,
    controlPi_85_4, controlPi_85_5, controlPi_85_6, controlPi_85_7,
    n2_ntk1, n11_ntk1, n13_ntk1, n16_ntk1, n21_ntk1, n45_ntk1, n46_ntk1,
    n55_ntk1, n74_ntk1, n75_ntk1, n81_ntk1, n84_ntk1, n85_ntk1, n93_ntk1,
    n96_ntk1, n98_ntk1, n101_ntk1, n111_ntk1, n128_ntk1, n131_ntk1,
    n134_ntk1, n139_ntk1, n153_ntk1, n159_ntk1, n177_ntk1, n199_ntk1,
    n206_ntk1, n211_ntk1, n216_ntk1, n223_ntk1, n243_ntk1, n264_ntk1,
    n266_ntk1, n280_ntk1, n282_ntk1, n287_ntk1, n290_ntk1, n309_ntk1,
    n336_ntk1, n346_ntk1, n349_ntk1, n360_ntk1, n368_ntk1, n369_ntk1,
    n377_ntk1, n388_ntk1, n394_ntk1, n409_ntk1, n428_ntk1, n435_ntk1,
    n447_ntk1, n454_ntk1, n457_ntk1, n468_ntk1, n471_ntk1, n481_ntk1,
    n494_ntk1, n500_ntk1, n507_ntk1, n511_ntk1, n519_ntk1, n525_ntk1,
    n557_ntk1, n561_ntk1, n569_ntk1, n571_ntk1, n575_ntk1, n581_ntk1,
    n582_ntk1, n583_ntk1, n587_ntk1, n600_ntk1, n603_ntk1, n609_ntk1,
    n613_ntk1, n614_ntk1, n616_ntk1, n646_ntk1, n659_ntk1, n661_ntk1,
    n664_ntk1, n673_ntk1;
  output miter;
  wire new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_,
    new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_,
    new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_,
    new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_,
    new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_,
    new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_,
    new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_,
    new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_,
    new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_,
    new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_,
    new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_,
    new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_,
    new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_,
    new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_,
    new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_,
    new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_,
    new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_,
    new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_,
    new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_,
    new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_,
    new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_,
    new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_,
    new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_,
    new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_,
    new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_,
    new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_,
    new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_,
    new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_,
    new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_,
    new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_,
    new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_,
    new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_,
    new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_,
    new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_,
    new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_,
    new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_,
    new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_,
    new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_,
    new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_,
    new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_,
    new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_,
    new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_,
    new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_,
    new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_,
    new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_,
    new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_,
    new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_,
    new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_,
    new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_,
    new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_,
    new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_,
    new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_,
    new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_,
    new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_,
    new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_,
    new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_,
    new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_,
    new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_,
    new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_,
    new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_,
    new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_,
    new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_,
    new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_,
    new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_,
    new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_,
    new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_,
    new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_,
    new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_,
    new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_,
    new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_,
    new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_,
    new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_,
    new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_,
    new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_,
    new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_,
    new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_,
    new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_,
    new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_,
    new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_,
    new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_,
    new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_,
    new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_,
    new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_,
    new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_,
    new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_,
    new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_,
    new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_,
    new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_,
    new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_,
    new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_,
    new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_,
    new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_,
    new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_,
    new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_,
    new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_,
    new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_,
    new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_,
    new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_,
    new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_,
    new_n1756_, new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_,
    new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_,
    new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_,
    new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_,
    new_n1780_, new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_,
    new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_,
    new_n1792_, new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_,
    new_n1798_, new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_,
    new_n1804_, new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_,
    new_n1810_, new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_,
    new_n1816_, new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_,
    new_n1822_, new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_,
    new_n1828_, new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_,
    new_n1834_, new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1839_,
    new_n1840_, new_n1841_, new_n1842_, new_n1843_, new_n1844_, new_n1845_,
    new_n1846_, new_n1847_, new_n1848_, new_n1849_, new_n1850_, new_n1851_,
    new_n1852_, new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_,
    new_n1858_, new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1863_,
    new_n1864_, new_n1865_, new_n1866_, new_n1867_, new_n1868_, new_n1869_,
    new_n1870_, new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_,
    new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1881_,
    new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1886_, new_n1887_,
    new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_,
    new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_,
    new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_,
    new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_,
    new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_,
    new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_,
    new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_, new_n1929_,
    new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_,
    new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_, new_n1941_,
    new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_,
    new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_, new_n1953_,
    new_n1954_, new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1959_,
    new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_,
    new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_,
    new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_,
    new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_,
    new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_,
    new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_,
    new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_,
    new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_,
    new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_,
    new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_,
    new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_,
    new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_,
    new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_,
    new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_,
    new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_,
    new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_,
    new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2061_,
    new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2067_,
    new_n2068_, new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_,
    new_n2074_, new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_,
    new_n2080_, new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2085_,
    new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_, new_n2091_,
    new_n2092_, new_n2093_, new_n2094_, new_n2095_, new_n2096_, new_n2097_,
    new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2102_, new_n2103_,
    new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_, new_n2109_,
    new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2115_,
    new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2121_,
    new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_,
    new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_,
    new_n2134_, new_n2135_, new_n2136_, new_n2137_, new_n2138_, new_n2139_,
    new_n2140_, new_n2141_, new_n2142_, new_n2143_, new_n2144_, new_n2145_,
    new_n2146_, new_n2147_, new_n2148_, new_n2149_, new_n2150_, new_n2151_,
    new_n2152_, new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_,
    new_n2158_, new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_,
    new_n2164_, new_n2165_, new_n2166_, new_n2167_, new_n2168_, new_n2169_,
    new_n2170_, new_n2171_, new_n2172_, new_n2173_, new_n2174_, new_n2175_,
    new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_,
    new_n2182_, new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_,
    new_n2188_, new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_,
    new_n2194_, new_n2195_, new_n2196_, new_n2197_, new_n2198_, new_n2199_,
    new_n2200_, new_n2201_, new_n2202_, new_n2203_, new_n2204_, new_n2205_,
    new_n2206_, new_n2207_, new_n2208_, new_n2209_, new_n2210_, new_n2211_,
    new_n2212_, new_n2213_, new_n2214_, new_n2215_, new_n2216_, new_n2217_,
    new_n2218_, new_n2219_, new_n2220_, new_n2221_, new_n2222_, new_n2223_,
    new_n2224_, new_n2225_, new_n2226_, new_n2227_, new_n2228_, new_n2229_,
    new_n2230_, new_n2231_, new_n2232_, new_n2233_, new_n2234_, new_n2235_,
    new_n2236_, new_n2237_, new_n2238_, new_n2239_, new_n2240_, new_n2241_,
    new_n2242_, new_n2243_, new_n2244_, new_n2245_, new_n2246_, new_n2247_,
    new_n2248_, new_n2249_, new_n2250_, new_n2251_, new_n2252_, new_n2253_,
    new_n2254_, new_n2255_, new_n2256_, new_n2257_, new_n2258_, new_n2259_,
    new_n2260_, new_n2261_, new_n2262_, new_n2263_, new_n2264_, new_n2265_,
    new_n2266_, new_n2267_, new_n2268_, new_n2269_, new_n2270_, new_n2271_,
    new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2276_, new_n2277_,
    new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_, new_n2283_,
    new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_, new_n2289_,
    new_n2290_, new_n2291_, new_n2292_, new_n2293_, new_n2294_, new_n2295_,
    new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_, new_n2301_,
    new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_, new_n2307_,
    new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_, new_n2313_,
    new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_, new_n2319_,
    new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_, new_n2325_,
    new_n2326_, new_n2327_, new_n2328_, new_n2329_, new_n2330_, new_n2331_,
    new_n2332_, new_n2333_, new_n2334_, new_n2335_, new_n2336_, new_n2337_,
    new_n2338_, new_n2339_, new_n2340_, new_n2341_, new_n2342_, new_n2343_,
    new_n2344_, new_n2345_, new_n2346_, new_n2347_, new_n2348_, new_n2349_,
    new_n2350_, new_n2351_, new_n2352_, new_n2353_, new_n2354_, new_n2355_,
    new_n2356_, new_n2357_, new_n2358_, new_n2359_, new_n2360_, new_n2361_,
    new_n2362_, new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_,
    new_n2368_, new_n2369_, new_n2370_, new_n2371_, new_n2372_, new_n2373_,
    new_n2374_, new_n2375_, new_n2376_, new_n2377_, new_n2378_, new_n2379_,
    new_n2380_, new_n2381_, new_n2382_, new_n2383_, new_n2384_, new_n2385_,
    new_n2386_, new_n2387_, new_n2388_, new_n2389_, new_n2390_, new_n2391_,
    new_n2392_, new_n2393_, new_n2394_, new_n2395_, new_n2396_, new_n2397_,
    new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_, new_n2403_,
    new_n2404_, new_n2405_, new_n2406_, new_n2407_, new_n2408_, new_n2409_,
    new_n2410_, new_n2411_, new_n2412_, new_n2413_, new_n2414_, new_n2415_,
    new_n2416_, new_n2417_, new_n2418_, new_n2419_, new_n2420_, new_n2421_,
    new_n2422_, new_n2423_, new_n2424_, new_n2425_, new_n2426_, new_n2427_,
    new_n2428_, new_n2429_, new_n2430_, new_n2431_, new_n2432_, new_n2433_,
    new_n2434_, new_n2435_, new_n2436_, new_n2437_, new_n2438_, new_n2439_,
    new_n2440_, new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_,
    new_n2446_, new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_,
    new_n2452_, new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_,
    new_n2458_, new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_,
    new_n2464_, new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_,
    new_n2470_, new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_,
    new_n2476_, new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_,
    new_n2482_, new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_,
    new_n2488_, new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_,
    new_n2494_, new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_,
    new_n2500_, new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_,
    new_n2506_, new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_,
    new_n2512_, new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_,
    new_n2518_, new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_,
    new_n2524_, new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_,
    new_n2530_, new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_,
    new_n2536_, new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_,
    new_n2542_, new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_,
    new_n2548_, new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_,
    new_n2554_, new_n2555_, new_n2556_, new_n2557_, new_n2558_, new_n2559_,
    new_n2560_, new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_,
    new_n2566_, new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_,
    new_n2572_, new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_,
    new_n2578_, new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_,
    new_n2584_, new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2589_,
    new_n2590_, new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_,
    new_n2596_, new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_,
    new_n2602_, new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_,
    new_n2608_, new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2613_,
    new_n2614_, new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2619_,
    new_n2620_, new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_,
    new_n2626_, new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_,
    new_n2632_, new_n2633_, new_n2634_, new_n2635_, new_n2636_, new_n2637_,
    new_n2638_, new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_,
    new_n2644_, new_n2645_, new_n2646_, new_n2647_, new_n2648_, new_n2649_,
    new_n2650_, new_n2651_, new_n2652_, new_n2653_, new_n2654_, new_n2655_,
    new_n2656_, new_n2657_, new_n2658_, new_n2659_, new_n2660_, new_n2661_,
    new_n2662_, new_n2663_, new_n2664_, new_n2665_, new_n2666_, new_n2667_,
    new_n2668_, new_n2669_, new_n2670_, new_n2671_, new_n2672_, new_n2673_,
    new_n2674_, new_n2675_, new_n2676_, new_n2677_, new_n2678_, new_n2679_,
    new_n2680_, new_n2681_, new_n2682_, new_n2683_, new_n2684_, new_n2685_,
    new_n2686_, new_n2687_, new_n2688_, new_n2689_, new_n2690_, new_n2691_,
    new_n2692_, new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_,
    new_n2698_, new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_,
    new_n2704_, new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2709_,
    new_n2710_, new_n2711_, new_n2712_, new_n2713_, new_n2714_, new_n2715_,
    new_n2716_, new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_,
    new_n2722_, new_n2723_, new_n2724_, new_n2725_, new_n2726_, new_n2727_,
    new_n2728_, new_n2729_, new_n2730_, new_n2731_, new_n2732_, new_n2733_,
    new_n2734_, new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_,
    new_n2740_, new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_,
    new_n2746_, new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_,
    new_n2752_, new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_,
    new_n2758_, new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2763_,
    new_n2764_, new_n2765_, new_n2766_, new_n2767_, new_n2768_, new_n2769_,
    new_n2770_, new_n2771_, new_n2772_, new_n2773_, new_n2774_, new_n2775_,
    new_n2776_, new_n2777_, new_n2778_, new_n2779_, new_n2780_, new_n2781_,
    new_n2782_, new_n2783_, new_n2784_, new_n2785_, new_n2786_, new_n2787_,
    new_n2788_, new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_,
    new_n2794_, new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_,
    new_n2800_, new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_,
    new_n2806_, new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_,
    new_n2812_, new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_,
    new_n2818_, new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2823_,
    new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_,
    new_n2830_, new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_,
    new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_,
    new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_,
    new_n2848_, new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_,
    new_n2854_, new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_,
    new_n2860_, new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_,
    new_n2866_, new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_,
    new_n2872_, new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_,
    new_n2878_, new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_,
    new_n2884_, new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_,
    new_n2890_, new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_,
    new_n2896_, new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_,
    new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2907_,
    new_n2908_, new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_,
    new_n2914_, new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_,
    new_n2920_, new_n2921_, new_n2922_, new_n2923_, new_n2924_, new_n2925_,
    new_n2926_, new_n2927_, new_n2928_, new_n2929_, new_n2930_, new_n2931_,
    new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2936_, new_n2937_,
    new_n2938_, new_n2939_, new_n2940_, new_n2941_, new_n2942_, new_n2943_,
    new_n2944_, new_n2945_, new_n2946_, new_n2947_, new_n2948_, new_n2949_,
    new_n2950_, new_n2951_, new_n2952_, new_n2953_, new_n2954_, new_n2955_,
    new_n2956_, new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2961_,
    new_n2962_, new_n2963_, new_n2964_, new_n2965_, new_n2966_, new_n2967_,
    new_n2968_, new_n2969_, new_n2970_, new_n2971_, new_n2972_, new_n2973_,
    new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_, new_n2979_,
    new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_, new_n2985_,
    new_n2986_, new_n2987_, new_n2988_, new_n2989_, new_n2990_, new_n2991_,
    new_n2992_, new_n2993_, new_n2994_, new_n2995_, new_n2996_, new_n2997_,
    new_n2998_, new_n2999_, new_n3000_, new_n3001_, new_n3002_, new_n3003_,
    new_n3004_, new_n3005_, new_n3006_, new_n3007_, new_n3008_, new_n3009_,
    new_n3010_, new_n3011_, new_n3012_, new_n3013_, new_n3014_, new_n3015_,
    new_n3016_, new_n3017_, new_n3018_, new_n3019_, new_n3020_, new_n3021_,
    new_n3022_, new_n3023_, new_n3024_, new_n3025_, new_n3026_, new_n3027_,
    new_n3028_, new_n3029_, new_n3030_, new_n3031_, new_n3032_, new_n3033_,
    new_n3034_, new_n3035_, new_n3036_, new_n3037_, new_n3038_, new_n3039_,
    new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3044_, new_n3045_,
    new_n3046_, new_n3047_, new_n3048_, new_n3049_, new_n3050_, new_n3051_,
    new_n3052_, new_n3053_, new_n3054_, new_n3055_, new_n3056_, new_n3057_,
    new_n3058_, new_n3059_, new_n3060_, new_n3061_, new_n3062_, new_n3063_,
    new_n3064_, new_n3065_, new_n3066_, new_n3067_, new_n3068_, new_n3069_,
    new_n3070_, new_n3071_, new_n3072_, new_n3073_, new_n3074_, new_n3075_,
    new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_, new_n3081_,
    new_n3082_, new_n3083_, new_n3084_, new_n3085_, new_n3086_, new_n3087_,
    new_n3088_, new_n3089_, new_n3090_, new_n3091_, new_n3092_, new_n3093_,
    new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3098_, new_n3099_,
    new_n3100_, new_n3101_, new_n3102_, new_n3103_, new_n3104_, new_n3105_,
    new_n3106_, new_n3107_, new_n3108_, new_n3109_, new_n3110_, new_n3111_,
    new_n3112_, new_n3113_, new_n3114_, new_n3115_, new_n3116_, new_n3117_,
    new_n3118_, new_n3119_, new_n3120_, new_n3121_, new_n3122_, new_n3123_,
    new_n3124_, new_n3125_, new_n3126_, new_n3127_, new_n3128_, new_n3129_,
    new_n3130_, new_n3131_, new_n3132_, new_n3133_, new_n3134_, new_n3135_,
    new_n3136_, new_n3137_, new_n3138_, new_n3139_, new_n3140_, new_n3141_,
    new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_, new_n3147_,
    new_n3148_, new_n3149_, new_n3150_, new_n3151_, new_n3152_, new_n3153_,
    new_n3154_, new_n3155_, new_n3156_, new_n3157_, new_n3158_, new_n3159_,
    new_n3160_, new_n3161_, new_n3162_, new_n3163_, new_n3164_, new_n3165_,
    new_n3166_, new_n3167_, new_n3168_, new_n3169_, new_n3170_, new_n3171_,
    new_n3172_, new_n3173_, new_n3174_, new_n3175_, new_n3176_, new_n3177_,
    new_n3178_, new_n3179_, new_n3180_, new_n3181_, new_n3182_, new_n3183_,
    new_n3184_, new_n3185_, new_n3186_, new_n3187_, new_n3188_, new_n3189_,
    new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_, new_n3195_,
    new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_, new_n3201_,
    new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_, new_n3207_,
    new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_, new_n3213_,
    new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_, new_n3219_,
    new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_, new_n3225_,
    new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_, new_n3231_,
    new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_, new_n3237_,
    new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_, new_n3243_,
    new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_, new_n3249_,
    new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_, new_n3255_,
    new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_, new_n3261_,
    new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_, new_n3267_,
    new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_, new_n3273_,
    new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_, new_n3279_,
    new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_, new_n3285_,
    new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_, new_n3291_,
    new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_, new_n3297_,
    new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_, new_n3303_,
    new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_, new_n3309_,
    new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_, new_n3315_,
    new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_, new_n3321_,
    new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_, new_n3327_,
    new_n3328_, new_n3329_, new_n3330_, new_n3331_, new_n3332_, new_n3333_,
    new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_, new_n3339_,
    new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_, new_n3345_,
    new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_, new_n3351_,
    new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_, new_n3357_,
    new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_, new_n3363_,
    new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_, new_n3369_,
    new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_, new_n3375_,
    new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_, new_n3381_,
    new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_, new_n3387_,
    new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_, new_n3393_,
    new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_, new_n3399_,
    new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_, new_n3405_,
    new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_, new_n3411_,
    new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_, new_n3417_,
    new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_,
    new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3428_, new_n3429_,
    new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3434_, new_n3435_,
    new_n3436_, new_n3437_, new_n3438_, new_n3439_, new_n3440_, new_n3441_,
    new_n3442_, new_n3443_, new_n3444_, new_n3445_, new_n3446_, new_n3447_,
    new_n3448_, new_n3449_, new_n3450_, new_n3451_, new_n3452_, new_n3453_,
    new_n3454_, new_n3455_, new_n3456_, new_n3457_, new_n3458_, new_n3459_,
    new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_, new_n3465_,
    new_n3466_, new_n3467_, new_n3468_, new_n3469_, new_n3470_, new_n3471_,
    new_n3472_, new_n3473_, new_n3474_, new_n3475_, new_n3476_, new_n3477_,
    new_n3478_, new_n3479_, new_n3480_, new_n3481_, new_n3482_, new_n3483_,
    new_n3484_, new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_,
    new_n3490_, new_n3491_, new_n3492_, new_n3493_, new_n3494_, new_n3495_,
    new_n3496_, new_n3497_, new_n3498_, new_n3499_, new_n3500_, new_n3501_,
    new_n3502_, new_n3503_, new_n3504_, new_n3505_, new_n3506_, new_n3507_,
    new_n3508_, new_n3509_, new_n3510_, new_n3511_, new_n3512_, new_n3513_,
    new_n3514_, new_n3515_, new_n3516_, new_n3517_, new_n3518_, new_n3519_,
    new_n3520_, new_n3521_, new_n3522_, new_n3523_, new_n3524_, new_n3525_,
    new_n3526_, new_n3527_, new_n3528_, new_n3529_, new_n3530_, new_n3531_,
    new_n3532_, new_n3533_, new_n3534_, new_n3535_, new_n3536_, new_n3537_,
    new_n3538_, new_n3539_, new_n3540_, new_n3541_, new_n3542_, new_n3543_,
    new_n3544_, new_n3545_, new_n3546_, new_n3547_, new_n3548_, new_n3549_,
    new_n3550_, new_n3551_, new_n3552_, new_n3553_, new_n3554_, new_n3555_,
    new_n3556_, new_n3557_, new_n3558_, new_n3559_, new_n3560_, new_n3561_,
    new_n3562_, new_n3563_, new_n3564_, new_n3565_, new_n3566_, new_n3567_,
    new_n3568_, new_n3569_, new_n3570_, new_n3571_, new_n3572_, new_n3573_,
    new_n3574_, new_n3575_, new_n3576_, new_n3577_, new_n3578_, new_n3579_,
    new_n3580_, new_n3581_, new_n3582_, new_n3583_, new_n3584_, new_n3585_,
    new_n3586_, new_n3587_, new_n3588_, new_n3589_, new_n3590_, new_n3591_,
    new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_, new_n3597_,
    new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3602_, new_n3603_,
    new_n3604_, new_n3605_, new_n3606_, new_n3607_, new_n3608_, new_n3609_,
    new_n3610_, new_n3611_, new_n3612_, new_n3613_, new_n3614_, new_n3615_,
    new_n3616_, new_n3617_, new_n3618_, new_n3619_, new_n3620_, new_n3621_,
    new_n3622_, new_n3623_, new_n3624_, new_n3625_, new_n3626_, new_n3627_,
    new_n3628_, new_n3629_, new_n3630_, new_n3631_, new_n3632_, new_n3633_,
    new_n3634_, new_n3635_, new_n3636_, new_n3637_, new_n3638_, new_n3639_,
    new_n3640_, new_n3641_, new_n3642_, new_n3643_, new_n3644_, new_n3645_,
    new_n3646_, new_n3647_, new_n3648_, new_n3649_, new_n3650_, new_n3651_,
    new_n3652_, new_n3653_, new_n3654_, new_n3655_, new_n3656_, new_n3657_,
    new_n3658_, new_n3659_, new_n3660_, new_n3661_, new_n3662_, new_n3663_,
    new_n3664_, new_n3665_, new_n3666_, new_n3667_, new_n3668_, new_n3669_,
    new_n3670_, new_n3671_, new_n3672_, new_n3673_, new_n3674_, new_n3675_,
    new_n3676_, new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3681_,
    new_n3682_, new_n3683_, new_n3684_, new_n3685_, new_n3686_, new_n3687_,
    new_n3688_, new_n3689_, new_n3690_, new_n3691_, new_n3692_, new_n3693_,
    new_n3694_, new_n3695_, new_n3696_, new_n3697_, new_n3698_, new_n3699_,
    new_n3700_, new_n3701_, new_n3702_, new_n3703_, new_n3704_, new_n3705_,
    new_n3706_, new_n3707_, new_n3708_, new_n3709_, new_n3710_, new_n3711_,
    new_n3712_, new_n3713_, new_n3714_, new_n3715_, new_n3716_, new_n3717_,
    new_n3718_, new_n3719_, new_n3720_, new_n3721_, new_n3722_, new_n3723_,
    new_n3724_, new_n3725_, new_n3726_, new_n3727_, new_n3728_, new_n3729_,
    new_n3730_, new_n3731_, new_n3732_, new_n3733_, new_n3734_, new_n3735_,
    new_n3736_, new_n3737_, new_n3738_, new_n3739_, new_n3740_, new_n3741_,
    new_n3742_, new_n3743_, new_n3744_, new_n3745_, new_n3746_, new_n3747_,
    new_n3748_, new_n3749_, new_n3750_, new_n3751_, new_n3752_, new_n3753_,
    new_n3754_, new_n3755_, new_n3756_, new_n3757_, new_n3758_, new_n3759_,
    new_n3760_, new_n3761_, new_n3762_, new_n3763_, new_n3764_, new_n3765_,
    new_n3766_, new_n3767_, new_n3768_, new_n3769_, new_n3770_, new_n3771_,
    new_n3772_, new_n3773_, new_n3774_, new_n3775_, new_n3776_, new_n3777_,
    new_n3778_, new_n3779_, new_n3780_, new_n3781_, new_n3782_, new_n3783_,
    new_n3784_, new_n3785_, new_n3786_, new_n3787_, new_n3788_, new_n3789_,
    new_n3790_, new_n3791_, new_n3792_, new_n3793_, new_n3794_, new_n3795_,
    new_n3796_, new_n3797_, new_n3798_, new_n3799_, new_n3800_, new_n3801_,
    new_n3802_, new_n3803_, new_n3804_, new_n3805_, new_n3806_, new_n3807_,
    new_n3808_, new_n3809_, new_n3810_, new_n3811_, new_n3812_, new_n3813_,
    new_n3814_, new_n3815_, new_n3816_, new_n3817_, new_n3818_, new_n3819_,
    new_n3820_, new_n3821_, new_n3822_, new_n3823_, new_n3824_, new_n3825_,
    new_n3826_, new_n3827_, new_n3828_, new_n3829_, new_n3830_, new_n3831_,
    new_n3832_, new_n3833_, new_n3834_, new_n3835_, new_n3836_, new_n3837_,
    new_n3838_, new_n3839_, new_n3840_, new_n3841_, new_n3842_, new_n3843_,
    new_n3844_, new_n3845_, new_n3846_, new_n3847_, new_n3848_, new_n3849_,
    new_n3850_, new_n3851_, new_n3852_, new_n3853_, new_n3854_, new_n3855_,
    new_n3856_, new_n3857_, new_n3858_, new_n3859_, new_n3860_, new_n3861_,
    new_n3862_, new_n3863_, new_n3864_, new_n3865_, new_n3866_, new_n3867_,
    new_n3868_, new_n3869_, new_n3870_, new_n3871_, new_n3872_, new_n3873_,
    new_n3874_, new_n3875_, new_n3876_, new_n3877_, new_n3878_, new_n3879_,
    new_n3880_, new_n3881_, new_n3882_, new_n3883_, new_n3884_, new_n3885_,
    new_n3886_, new_n3887_, new_n3888_, new_n3889_, new_n3890_, new_n3891_,
    new_n3892_, new_n3893_, new_n3894_, new_n3895_, new_n3896_, new_n3897_,
    new_n3898_, new_n3899_, new_n3900_, new_n3901_, new_n3902_, new_n3903_,
    new_n3904_, new_n3905_, new_n3906_, new_n3907_, new_n3908_, new_n3909_,
    new_n3910_, new_n3911_, new_n3912_, new_n3913_, new_n3914_, new_n3915_,
    new_n3916_, new_n3917_, new_n3918_, new_n3919_, new_n3920_, new_n3921_,
    new_n3922_, new_n3923_, new_n3924_, new_n3925_, new_n3926_, new_n3927_,
    new_n3928_, new_n3929_, new_n3930_, new_n3931_, new_n3932_, new_n3933_,
    new_n3934_, new_n3935_, new_n3936_, new_n3937_, new_n3938_, new_n3939_,
    new_n3940_, new_n3941_, new_n3942_, new_n3943_, new_n3944_, new_n3945_,
    new_n3946_, new_n3947_, new_n3948_, new_n3949_, new_n3950_, new_n3951_,
    new_n3952_, new_n3953_, new_n3954_, new_n3955_, new_n3956_, new_n3957_,
    new_n3958_, new_n3959_, new_n3960_, new_n3961_, new_n3962_, new_n3963_,
    new_n3964_, new_n3965_, new_n3966_, new_n3967_, new_n3968_, new_n3969_,
    new_n3970_, new_n3971_, new_n3972_, new_n3973_, new_n3974_, new_n3975_;
  assign new_n772_ = ~n206_ntk1 & ~n368_ntk1;
  assign new_n773_ = n2_ntk1 & n582_ntk1;
  assign new_n774_ = n287_ntk1 & n600_ntk1;
  assign new_n775_ = ~n2_ntk1 & ~n582_ntk1;
  assign new_n776_ = new_n774_ & ~new_n775_;
  assign new_n777_ = ~new_n773_ & ~new_n776_;
  assign new_n778_ = ~n75_ntk1 & ~n435_ntk1;
  assign new_n779_ = n75_ntk1 & n435_ntk1;
  assign new_n780_ = ~new_n778_ & ~new_n779_;
  assign new_n781_ = new_n777_ & ~new_n780_;
  assign new_n782_ = ~new_n777_ & new_n780_;
  assign new_n783_ = n349_ntk1 & ~new_n782_;
  assign new_n784_ = ~new_n781_ & new_n783_;
  assign new_n785_ = n2_ntk1 & n13_ntk1;
  assign new_n786_ = n280_ntk1 & n287_ntk1;
  assign new_n787_ = ~n2_ntk1 & ~n13_ntk1;
  assign new_n788_ = new_n786_ & ~new_n787_;
  assign new_n789_ = ~new_n785_ & ~new_n788_;
  assign new_n790_ = ~n75_ntk1 & ~n177_ntk1;
  assign new_n791_ = n75_ntk1 & n177_ntk1;
  assign new_n792_ = ~new_n790_ & ~new_n791_;
  assign new_n793_ = ~new_n789_ & new_n792_;
  assign new_n794_ = n85_ntk1 & ~n349_ntk1;
  assign new_n795_ = new_n789_ & ~new_n792_;
  assign new_n796_ = new_n794_ & ~new_n795_;
  assign new_n797_ = ~new_n793_ & new_n796_;
  assign new_n798_ = ~n85_ntk1 & ~n349_ntk1;
  assign new_n799_ = n211_ntk1 & new_n798_;
  assign new_n800_ = ~new_n797_ & ~new_n799_;
  assign new_n801_ = ~new_n784_ & new_n800_;
  assign new_n802_ = new_n772_ & ~new_n801_;
  assign new_n803_ = n454_ntk1 & n659_ntk1;
  assign new_n804_ = ~n216_ntk1 & ~new_n803_;
  assign new_n805_ = n216_ntk1 & new_n803_;
  assign new_n806_ = ~new_n804_ & ~new_n805_;
  assign new_n807_ = n206_ntk1 & new_n806_;
  assign new_n808_ = n2_ntk1 & n159_ntk1;
  assign new_n809_ = n96_ntk1 & n287_ntk1;
  assign new_n810_ = ~n2_ntk1 & ~n159_ntk1;
  assign new_n811_ = new_n809_ & ~new_n810_;
  assign new_n812_ = ~new_n808_ & ~new_n811_;
  assign new_n813_ = ~n75_ntk1 & ~n131_ntk1;
  assign new_n814_ = n75_ntk1 & n131_ntk1;
  assign new_n815_ = ~new_n813_ & ~new_n814_;
  assign new_n816_ = new_n812_ & ~new_n815_;
  assign new_n817_ = ~n206_ntk1 & n368_ntk1;
  assign new_n818_ = ~new_n812_ & new_n815_;
  assign new_n819_ = new_n817_ & ~new_n818_;
  assign new_n820_ = ~new_n816_ & new_n819_;
  assign new_n821_ = ~new_n807_ & ~new_n820_;
  assign new_n822_ = ~new_n802_ & new_n821_;
  assign new_n823_ = ~n93_ntk1 & ~new_n822_;
  assign new_n824_ = n428_ntk1 & n454_ntk1;
  assign new_n825_ = n409_ntk1 & ~n428_ntk1;
  assign new_n826_ = ~n409_ntk1 & n428_ntk1;
  assign new_n827_ = ~new_n825_ & ~new_n826_;
  assign new_n828_ = n216_ntk1 & ~new_n827_;
  assign new_n829_ = ~n216_ntk1 & new_n827_;
  assign new_n830_ = ~new_n828_ & ~new_n829_;
  assign new_n831_ = ~new_n824_ & ~new_n830_;
  assign new_n832_ = new_n824_ & new_n830_;
  assign new_n833_ = ~new_n831_ & ~new_n832_;
  assign new_n834_ = n93_ntk1 & new_n833_;
  assign new_n835_ = ~new_n823_ & ~new_n834_;
  assign new_n836_ = n511_ntk1 & ~n659_ntk1;
  assign new_n837_ = ~n454_ntk1 & new_n836_;
  assign new_n838_ = n216_ntk1 & ~new_n837_;
  assign new_n839_ = ~n216_ntk1 & new_n837_;
  assign new_n840_ = ~new_n838_ & ~new_n839_;
  assign new_n841_ = n266_ntk1 & new_n840_;
  assign new_n842_ = ~n266_ntk1 & ~n457_ntk1;
  assign new_n843_ = ~new_n841_ & ~new_n842_;
  assign new_n844_ = ~new_n835_ & ~new_n843_;
  assign new_n845_ = new_n835_ & new_n843_;
  assign new_n846_ = ~new_n844_ & ~new_n845_;
  assign new_n847_ = n93_ntk1 & n659_ntk1;
  assign new_n848_ = ~n280_ntk1 & ~n287_ntk1;
  assign new_n849_ = ~new_n786_ & ~new_n848_;
  assign new_n850_ = new_n794_ & new_n849_;
  assign new_n851_ = n664_ntk1 & new_n798_;
  assign new_n852_ = ~n287_ntk1 & ~n600_ntk1;
  assign new_n853_ = ~new_n774_ & ~new_n852_;
  assign new_n854_ = n349_ntk1 & new_n853_;
  assign new_n855_ = ~new_n851_ & ~new_n854_;
  assign new_n856_ = ~new_n850_ & new_n855_;
  assign new_n857_ = new_n772_ & ~new_n856_;
  assign new_n858_ = n206_ntk1 & ~n659_ntk1;
  assign new_n859_ = ~n96_ntk1 & ~n287_ntk1;
  assign new_n860_ = ~new_n809_ & new_n817_;
  assign new_n861_ = ~new_n859_ & new_n860_;
  assign new_n862_ = ~new_n858_ & ~new_n861_;
  assign new_n863_ = ~new_n857_ & new_n862_;
  assign new_n864_ = ~n93_ntk1 & ~new_n863_;
  assign new_n865_ = ~new_n847_ & ~new_n864_;
  assign new_n866_ = ~n511_ntk1 & n659_ntk1;
  assign new_n867_ = ~new_n836_ & ~new_n866_;
  assign new_n868_ = n266_ntk1 & ~new_n867_;
  assign new_n869_ = ~n266_ntk1 & n673_ntk1;
  assign new_n870_ = ~new_n868_ & ~new_n869_;
  assign new_n871_ = ~new_n865_ & new_n870_;
  assign new_n872_ = ~n428_ntk1 & ~n454_ntk1;
  assign new_n873_ = ~new_n824_ & ~new_n872_;
  assign new_n874_ = n93_ntk1 & new_n873_;
  assign new_n875_ = ~new_n785_ & ~new_n787_;
  assign new_n876_ = new_n786_ & ~new_n875_;
  assign new_n877_ = ~new_n786_ & new_n875_;
  assign new_n878_ = ~new_n876_ & ~new_n877_;
  assign new_n879_ = new_n794_ & ~new_n878_;
  assign new_n880_ = ~new_n773_ & ~new_n775_;
  assign new_n881_ = new_n774_ & ~new_n880_;
  assign new_n882_ = ~new_n774_ & new_n880_;
  assign new_n883_ = ~new_n881_ & ~new_n882_;
  assign new_n884_ = n349_ntk1 & ~new_n883_;
  assign new_n885_ = n525_ntk1 & new_n798_;
  assign new_n886_ = ~new_n884_ & ~new_n885_;
  assign new_n887_ = ~new_n879_ & new_n886_;
  assign new_n888_ = new_n772_ & ~new_n887_;
  assign new_n889_ = ~new_n808_ & ~new_n810_;
  assign new_n890_ = new_n809_ & ~new_n889_;
  assign new_n891_ = ~new_n809_ & new_n889_;
  assign new_n892_ = ~new_n890_ & ~new_n891_;
  assign new_n893_ = new_n817_ & ~new_n892_;
  assign new_n894_ = ~n454_ntk1 & ~n659_ntk1;
  assign new_n895_ = n206_ntk1 & ~new_n803_;
  assign new_n896_ = ~new_n894_ & new_n895_;
  assign new_n897_ = ~new_n893_ & ~new_n896_;
  assign new_n898_ = ~new_n888_ & new_n897_;
  assign new_n899_ = ~n93_ntk1 & ~new_n898_;
  assign new_n900_ = ~new_n874_ & ~new_n899_;
  assign new_n901_ = n454_ntk1 & ~new_n836_;
  assign new_n902_ = ~new_n837_ & ~new_n901_;
  assign new_n903_ = n266_ntk1 & new_n902_;
  assign new_n904_ = ~n46_ntk1 & ~n266_ntk1;
  assign new_n905_ = ~new_n903_ & ~new_n904_;
  assign new_n906_ = ~new_n900_ & ~new_n905_;
  assign new_n907_ = ~new_n871_ & ~new_n906_;
  assign new_n908_ = new_n900_ & new_n905_;
  assign new_n909_ = ~new_n907_ & ~new_n908_;
  assign new_n910_ = n266_ntk1 & new_n909_;
  assign new_n911_ = ~new_n900_ & new_n905_;
  assign new_n912_ = new_n900_ & ~new_n905_;
  assign new_n913_ = ~new_n865_ & ~new_n870_;
  assign new_n914_ = ~new_n912_ & new_n913_;
  assign new_n915_ = ~new_n911_ & ~new_n914_;
  assign new_n916_ = ~n266_ntk1 & ~new_n915_;
  assign new_n917_ = ~new_n910_ & ~new_n916_;
  assign new_n918_ = new_n846_ & new_n917_;
  assign new_n919_ = ~new_n846_ & ~new_n917_;
  assign new_n920_ = ~new_n918_ & ~new_n919_;
  assign new_n921_ = ~controlPi_69_1 & ~n349_ntk1;
  assign new_n922_ = controlPi_69_1 & ~n368_ntk1;
  assign new_n923_ = ~new_n921_ & ~new_n922_;
  assign new_n924_ = controlPi_69_3 & ~new_n923_;
  assign new_n925_ = ~controlPi_69_1 & ~n85_ntk1;
  assign new_n926_ = controlPi_69_1 & ~n93_ntk1;
  assign new_n927_ = ~new_n925_ & ~new_n926_;
  assign new_n928_ = ~controlPi_69_3 & ~new_n927_;
  assign new_n929_ = ~new_n924_ & ~new_n928_;
  assign new_n930_ = ~controlPi_69_2 & ~new_n929_;
  assign new_n931_ = ~controlPi_69_1 & ~n206_ntk1;
  assign new_n932_ = controlPi_69_1 & ~n266_ntk1;
  assign new_n933_ = ~new_n931_ & ~new_n932_;
  assign new_n934_ = controlPi_69_2 & ~new_n933_;
  assign new_n935_ = ~controlPi_69_3 & new_n934_;
  assign new_n936_ = ~new_n930_ & ~new_n935_;
  assign new_n937_ = controlPi_69_0 & ~new_n936_;
  assign new_n938_ = ~controlPi_69_0 & new_n936_;
  assign new_n939_ = ~new_n937_ & ~new_n938_;
  assign new_n940_ = ~controlPi_77_1 & ~n199_ntk1;
  assign new_n941_ = controlPi_77_1 & ~n211_ntk1;
  assign new_n942_ = ~new_n940_ & ~new_n941_;
  assign new_n943_ = ~controlPi_77_2 & new_n942_;
  assign new_n944_ = ~controlPi_77_1 & ~n216_ntk1;
  assign new_n945_ = controlPi_77_1 & ~n280_ntk1;
  assign new_n946_ = ~new_n944_ & ~new_n945_;
  assign new_n947_ = controlPi_77_2 & new_n946_;
  assign new_n948_ = ~new_n943_ & ~new_n947_;
  assign new_n949_ = ~controlPi_77_3 & new_n948_;
  assign new_n950_ = ~controlPi_77_1 & ~n287_ntk1;
  assign new_n951_ = controlPi_77_1 & ~n409_ntk1;
  assign new_n952_ = ~new_n950_ & ~new_n951_;
  assign new_n953_ = ~controlPi_77_2 & new_n952_;
  assign new_n954_ = ~controlPi_77_1 & ~n428_ntk1;
  assign new_n955_ = controlPi_77_1 & ~n435_ntk1;
  assign new_n956_ = ~new_n954_ & ~new_n955_;
  assign new_n957_ = controlPi_77_2 & new_n956_;
  assign new_n958_ = ~new_n953_ & ~new_n957_;
  assign new_n959_ = controlPi_77_3 & new_n958_;
  assign new_n960_ = ~new_n949_ & ~new_n959_;
  assign new_n961_ = controlPi_77_4 & ~new_n960_;
  assign new_n962_ = ~controlPi_77_1 & ~n2_ntk1;
  assign new_n963_ = controlPi_77_1 & ~n13_ntk1;
  assign new_n964_ = ~new_n962_ & ~new_n963_;
  assign new_n965_ = ~controlPi_77_2 & new_n964_;
  assign new_n966_ = ~controlPi_77_1 & ~n46_ntk1;
  assign new_n967_ = controlPi_77_1 & ~n75_ntk1;
  assign new_n968_ = ~new_n966_ & ~new_n967_;
  assign new_n969_ = controlPi_77_2 & new_n968_;
  assign new_n970_ = ~new_n965_ & ~new_n969_;
  assign new_n971_ = ~controlPi_77_3 & new_n970_;
  assign new_n972_ = ~controlPi_77_1 & ~n96_ntk1;
  assign new_n973_ = controlPi_77_1 & ~n131_ntk1;
  assign new_n974_ = ~new_n972_ & ~new_n973_;
  assign new_n975_ = ~controlPi_77_2 & new_n974_;
  assign new_n976_ = ~controlPi_77_1 & ~n159_ntk1;
  assign new_n977_ = controlPi_77_1 & ~n177_ntk1;
  assign new_n978_ = ~new_n976_ & ~new_n977_;
  assign new_n979_ = controlPi_77_2 & new_n978_;
  assign new_n980_ = ~new_n975_ & ~new_n979_;
  assign new_n981_ = controlPi_77_3 & new_n980_;
  assign new_n982_ = ~new_n971_ & ~new_n981_;
  assign new_n983_ = ~controlPi_77_4 & ~new_n982_;
  assign new_n984_ = ~new_n961_ & ~new_n983_;
  assign new_n985_ = ~controlPi_77_5 & ~new_n984_;
  assign new_n986_ = controlPi_77_1 & n659_ntk1;
  assign new_n987_ = ~controlPi_77_1 & n616_ntk1;
  assign new_n988_ = ~new_n986_ & ~new_n987_;
  assign new_n989_ = ~controlPi_77_2 & new_n988_;
  assign new_n990_ = controlPi_77_1 & n673_ntk1;
  assign new_n991_ = ~controlPi_77_1 & n664_ntk1;
  assign new_n992_ = ~new_n990_ & ~new_n991_;
  assign new_n993_ = controlPi_77_2 & new_n992_;
  assign new_n994_ = ~new_n989_ & ~new_n993_;
  assign new_n995_ = controlPi_77_4 & ~new_n994_;
  assign new_n996_ = controlPi_77_1 & n457_ntk1;
  assign new_n997_ = ~controlPi_77_1 & n454_ntk1;
  assign new_n998_ = ~new_n996_ & ~new_n997_;
  assign new_n999_ = ~controlPi_77_2 & new_n998_;
  assign new_n1000_ = controlPi_77_1 & n507_ntk1;
  assign new_n1001_ = ~controlPi_77_1 & n468_ntk1;
  assign new_n1002_ = ~new_n1000_ & ~new_n1001_;
  assign new_n1003_ = controlPi_77_2 & new_n1002_;
  assign new_n1004_ = ~new_n999_ & ~new_n1003_;
  assign new_n1005_ = ~controlPi_77_4 & ~new_n1004_;
  assign new_n1006_ = ~new_n995_ & ~new_n1005_;
  assign new_n1007_ = ~controlPi_77_3 & ~new_n1006_;
  assign new_n1008_ = controlPi_77_1 & n600_ntk1;
  assign new_n1009_ = ~controlPi_77_1 & n582_ntk1;
  assign new_n1010_ = ~new_n1008_ & ~new_n1009_;
  assign new_n1011_ = controlPi_77_2 & new_n1010_;
  assign new_n1012_ = controlPi_77_1 & n525_ntk1;
  assign new_n1013_ = ~controlPi_77_1 & n511_ntk1;
  assign new_n1014_ = ~new_n1012_ & ~new_n1013_;
  assign new_n1015_ = ~controlPi_77_2 & new_n1014_;
  assign new_n1016_ = ~new_n1011_ & ~new_n1015_;
  assign new_n1017_ = controlPi_77_3 & ~new_n1016_;
  assign new_n1018_ = ~controlPi_77_4 & new_n1017_;
  assign new_n1019_ = ~new_n1007_ & ~new_n1018_;
  assign new_n1020_ = controlPi_77_5 & ~new_n1019_;
  assign new_n1021_ = ~new_n985_ & ~new_n1020_;
  assign new_n1022_ = controlPi_77_0 & ~new_n1021_;
  assign new_n1023_ = ~controlPi_77_0 & new_n1021_;
  assign new_n1024_ = ~new_n1022_ & ~new_n1023_;
  assign new_n1025_ = new_n939_ & ~new_n1024_;
  assign new_n1026_ = ~controlPi_0_1 & ~n199_ntk1;
  assign new_n1027_ = controlPi_0_1 & ~n211_ntk1;
  assign new_n1028_ = ~new_n1026_ & ~new_n1027_;
  assign new_n1029_ = ~controlPi_0_2 & new_n1028_;
  assign new_n1030_ = ~controlPi_0_1 & ~n216_ntk1;
  assign new_n1031_ = controlPi_0_1 & ~n280_ntk1;
  assign new_n1032_ = ~new_n1030_ & ~new_n1031_;
  assign new_n1033_ = controlPi_0_2 & new_n1032_;
  assign new_n1034_ = ~new_n1029_ & ~new_n1033_;
  assign new_n1035_ = ~controlPi_0_3 & new_n1034_;
  assign new_n1036_ = ~controlPi_0_1 & ~n287_ntk1;
  assign new_n1037_ = controlPi_0_1 & ~n409_ntk1;
  assign new_n1038_ = ~new_n1036_ & ~new_n1037_;
  assign new_n1039_ = ~controlPi_0_2 & new_n1038_;
  assign new_n1040_ = ~controlPi_0_1 & ~n428_ntk1;
  assign new_n1041_ = controlPi_0_1 & ~n435_ntk1;
  assign new_n1042_ = ~new_n1040_ & ~new_n1041_;
  assign new_n1043_ = controlPi_0_2 & new_n1042_;
  assign new_n1044_ = ~new_n1039_ & ~new_n1043_;
  assign new_n1045_ = controlPi_0_3 & new_n1044_;
  assign new_n1046_ = ~new_n1035_ & ~new_n1045_;
  assign new_n1047_ = controlPi_0_4 & ~new_n1046_;
  assign new_n1048_ = ~controlPi_0_1 & ~n2_ntk1;
  assign new_n1049_ = controlPi_0_1 & ~n13_ntk1;
  assign new_n1050_ = ~new_n1048_ & ~new_n1049_;
  assign new_n1051_ = ~controlPi_0_2 & new_n1050_;
  assign new_n1052_ = ~controlPi_0_1 & ~n46_ntk1;
  assign new_n1053_ = controlPi_0_1 & ~n75_ntk1;
  assign new_n1054_ = ~new_n1052_ & ~new_n1053_;
  assign new_n1055_ = controlPi_0_2 & new_n1054_;
  assign new_n1056_ = ~new_n1051_ & ~new_n1055_;
  assign new_n1057_ = ~controlPi_0_3 & new_n1056_;
  assign new_n1058_ = ~controlPi_0_1 & ~n96_ntk1;
  assign new_n1059_ = controlPi_0_1 & ~n131_ntk1;
  assign new_n1060_ = ~new_n1058_ & ~new_n1059_;
  assign new_n1061_ = ~controlPi_0_2 & new_n1060_;
  assign new_n1062_ = ~controlPi_0_1 & ~n159_ntk1;
  assign new_n1063_ = controlPi_0_1 & ~n177_ntk1;
  assign new_n1064_ = ~new_n1062_ & ~new_n1063_;
  assign new_n1065_ = controlPi_0_2 & new_n1064_;
  assign new_n1066_ = ~new_n1061_ & ~new_n1065_;
  assign new_n1067_ = controlPi_0_3 & new_n1066_;
  assign new_n1068_ = ~new_n1057_ & ~new_n1067_;
  assign new_n1069_ = ~controlPi_0_4 & ~new_n1068_;
  assign new_n1070_ = ~new_n1047_ & ~new_n1069_;
  assign new_n1071_ = ~controlPi_0_5 & ~new_n1070_;
  assign new_n1072_ = controlPi_0_1 & n659_ntk1;
  assign new_n1073_ = ~controlPi_0_1 & n616_ntk1;
  assign new_n1074_ = ~new_n1072_ & ~new_n1073_;
  assign new_n1075_ = ~controlPi_0_2 & new_n1074_;
  assign new_n1076_ = controlPi_0_1 & n673_ntk1;
  assign new_n1077_ = ~controlPi_0_1 & n664_ntk1;
  assign new_n1078_ = ~new_n1076_ & ~new_n1077_;
  assign new_n1079_ = controlPi_0_2 & new_n1078_;
  assign new_n1080_ = ~new_n1075_ & ~new_n1079_;
  assign new_n1081_ = controlPi_0_4 & ~new_n1080_;
  assign new_n1082_ = controlPi_0_1 & n457_ntk1;
  assign new_n1083_ = ~controlPi_0_1 & n454_ntk1;
  assign new_n1084_ = ~new_n1082_ & ~new_n1083_;
  assign new_n1085_ = ~controlPi_0_2 & new_n1084_;
  assign new_n1086_ = controlPi_0_1 & n507_ntk1;
  assign new_n1087_ = ~controlPi_0_1 & n468_ntk1;
  assign new_n1088_ = ~new_n1086_ & ~new_n1087_;
  assign new_n1089_ = controlPi_0_2 & new_n1088_;
  assign new_n1090_ = ~new_n1085_ & ~new_n1089_;
  assign new_n1091_ = ~controlPi_0_4 & ~new_n1090_;
  assign new_n1092_ = ~new_n1081_ & ~new_n1091_;
  assign new_n1093_ = ~controlPi_0_3 & ~new_n1092_;
  assign new_n1094_ = controlPi_0_1 & n600_ntk1;
  assign new_n1095_ = ~controlPi_0_1 & n582_ntk1;
  assign new_n1096_ = ~new_n1094_ & ~new_n1095_;
  assign new_n1097_ = controlPi_0_2 & new_n1096_;
  assign new_n1098_ = controlPi_0_1 & n525_ntk1;
  assign new_n1099_ = ~controlPi_0_1 & n511_ntk1;
  assign new_n1100_ = ~new_n1098_ & ~new_n1099_;
  assign new_n1101_ = ~controlPi_0_2 & new_n1100_;
  assign new_n1102_ = ~new_n1097_ & ~new_n1101_;
  assign new_n1103_ = controlPi_0_3 & ~new_n1102_;
  assign new_n1104_ = ~controlPi_0_4 & new_n1103_;
  assign new_n1105_ = ~new_n1093_ & ~new_n1104_;
  assign new_n1106_ = controlPi_0_5 & ~new_n1105_;
  assign new_n1107_ = ~new_n1071_ & ~new_n1106_;
  assign new_n1108_ = controlPi_0_0 & ~new_n1107_;
  assign new_n1109_ = ~controlPi_0_0 & new_n1107_;
  assign new_n1110_ = ~new_n1108_ & ~new_n1109_;
  assign new_n1111_ = ~controlPi_70_1 & ~n199_ntk1;
  assign new_n1112_ = controlPi_70_1 & ~n211_ntk1;
  assign new_n1113_ = ~new_n1111_ & ~new_n1112_;
  assign new_n1114_ = ~controlPi_70_2 & new_n1113_;
  assign new_n1115_ = ~controlPi_70_1 & ~n216_ntk1;
  assign new_n1116_ = controlPi_70_1 & ~n280_ntk1;
  assign new_n1117_ = ~new_n1115_ & ~new_n1116_;
  assign new_n1118_ = controlPi_70_2 & new_n1117_;
  assign new_n1119_ = ~new_n1114_ & ~new_n1118_;
  assign new_n1120_ = ~controlPi_70_3 & new_n1119_;
  assign new_n1121_ = ~controlPi_70_1 & ~n287_ntk1;
  assign new_n1122_ = controlPi_70_1 & ~n409_ntk1;
  assign new_n1123_ = ~new_n1121_ & ~new_n1122_;
  assign new_n1124_ = ~controlPi_70_2 & new_n1123_;
  assign new_n1125_ = ~controlPi_70_1 & ~n428_ntk1;
  assign new_n1126_ = controlPi_70_1 & ~n435_ntk1;
  assign new_n1127_ = ~new_n1125_ & ~new_n1126_;
  assign new_n1128_ = controlPi_70_2 & new_n1127_;
  assign new_n1129_ = ~new_n1124_ & ~new_n1128_;
  assign new_n1130_ = controlPi_70_3 & new_n1129_;
  assign new_n1131_ = ~new_n1120_ & ~new_n1130_;
  assign new_n1132_ = controlPi_70_4 & ~new_n1131_;
  assign new_n1133_ = ~controlPi_70_1 & ~n2_ntk1;
  assign new_n1134_ = controlPi_70_1 & ~n13_ntk1;
  assign new_n1135_ = ~new_n1133_ & ~new_n1134_;
  assign new_n1136_ = ~controlPi_70_2 & new_n1135_;
  assign new_n1137_ = ~controlPi_70_1 & ~n46_ntk1;
  assign new_n1138_ = controlPi_70_1 & ~n75_ntk1;
  assign new_n1139_ = ~new_n1137_ & ~new_n1138_;
  assign new_n1140_ = controlPi_70_2 & new_n1139_;
  assign new_n1141_ = ~new_n1136_ & ~new_n1140_;
  assign new_n1142_ = ~controlPi_70_3 & new_n1141_;
  assign new_n1143_ = ~controlPi_70_1 & ~n96_ntk1;
  assign new_n1144_ = controlPi_70_1 & ~n131_ntk1;
  assign new_n1145_ = ~new_n1143_ & ~new_n1144_;
  assign new_n1146_ = ~controlPi_70_2 & new_n1145_;
  assign new_n1147_ = ~controlPi_70_1 & ~n159_ntk1;
  assign new_n1148_ = controlPi_70_1 & ~n177_ntk1;
  assign new_n1149_ = ~new_n1147_ & ~new_n1148_;
  assign new_n1150_ = controlPi_70_2 & new_n1149_;
  assign new_n1151_ = ~new_n1146_ & ~new_n1150_;
  assign new_n1152_ = controlPi_70_3 & new_n1151_;
  assign new_n1153_ = ~new_n1142_ & ~new_n1152_;
  assign new_n1154_ = ~controlPi_70_4 & ~new_n1153_;
  assign new_n1155_ = ~new_n1132_ & ~new_n1154_;
  assign new_n1156_ = ~controlPi_70_5 & ~new_n1155_;
  assign new_n1157_ = controlPi_70_1 & n659_ntk1;
  assign new_n1158_ = ~controlPi_70_1 & n616_ntk1;
  assign new_n1159_ = ~new_n1157_ & ~new_n1158_;
  assign new_n1160_ = ~controlPi_70_2 & new_n1159_;
  assign new_n1161_ = controlPi_70_1 & n673_ntk1;
  assign new_n1162_ = ~controlPi_70_1 & n664_ntk1;
  assign new_n1163_ = ~new_n1161_ & ~new_n1162_;
  assign new_n1164_ = controlPi_70_2 & new_n1163_;
  assign new_n1165_ = ~new_n1160_ & ~new_n1164_;
  assign new_n1166_ = controlPi_70_4 & ~new_n1165_;
  assign new_n1167_ = controlPi_70_1 & n457_ntk1;
  assign new_n1168_ = ~controlPi_70_1 & n454_ntk1;
  assign new_n1169_ = ~new_n1167_ & ~new_n1168_;
  assign new_n1170_ = ~controlPi_70_2 & new_n1169_;
  assign new_n1171_ = controlPi_70_1 & n507_ntk1;
  assign new_n1172_ = ~controlPi_70_1 & n468_ntk1;
  assign new_n1173_ = ~new_n1171_ & ~new_n1172_;
  assign new_n1174_ = controlPi_70_2 & new_n1173_;
  assign new_n1175_ = ~new_n1170_ & ~new_n1174_;
  assign new_n1176_ = ~controlPi_70_4 & ~new_n1175_;
  assign new_n1177_ = ~new_n1166_ & ~new_n1176_;
  assign new_n1178_ = ~controlPi_70_3 & ~new_n1177_;
  assign new_n1179_ = controlPi_70_1 & n600_ntk1;
  assign new_n1180_ = ~controlPi_70_1 & n582_ntk1;
  assign new_n1181_ = ~new_n1179_ & ~new_n1180_;
  assign new_n1182_ = controlPi_70_2 & new_n1181_;
  assign new_n1183_ = controlPi_70_1 & n525_ntk1;
  assign new_n1184_ = ~controlPi_70_1 & n511_ntk1;
  assign new_n1185_ = ~new_n1183_ & ~new_n1184_;
  assign new_n1186_ = ~controlPi_70_2 & new_n1185_;
  assign new_n1187_ = ~new_n1182_ & ~new_n1186_;
  assign new_n1188_ = controlPi_70_3 & ~new_n1187_;
  assign new_n1189_ = ~controlPi_70_4 & new_n1188_;
  assign new_n1190_ = ~new_n1178_ & ~new_n1189_;
  assign new_n1191_ = controlPi_70_5 & ~new_n1190_;
  assign new_n1192_ = ~new_n1156_ & ~new_n1191_;
  assign new_n1193_ = controlPi_70_0 & ~new_n1192_;
  assign new_n1194_ = ~controlPi_70_0 & new_n1192_;
  assign new_n1195_ = ~new_n1193_ & ~new_n1194_;
  assign new_n1196_ = ~new_n1110_ & ~new_n1195_;
  assign new_n1197_ = ~controlPi_17_1 & ~n199_ntk1;
  assign new_n1198_ = controlPi_17_1 & ~n211_ntk1;
  assign new_n1199_ = ~new_n1197_ & ~new_n1198_;
  assign new_n1200_ = ~controlPi_17_2 & new_n1199_;
  assign new_n1201_ = ~controlPi_17_1 & ~n216_ntk1;
  assign new_n1202_ = controlPi_17_1 & ~n280_ntk1;
  assign new_n1203_ = ~new_n1201_ & ~new_n1202_;
  assign new_n1204_ = controlPi_17_2 & new_n1203_;
  assign new_n1205_ = ~new_n1200_ & ~new_n1204_;
  assign new_n1206_ = ~controlPi_17_3 & new_n1205_;
  assign new_n1207_ = ~controlPi_17_1 & ~n287_ntk1;
  assign new_n1208_ = controlPi_17_1 & ~n409_ntk1;
  assign new_n1209_ = ~new_n1207_ & ~new_n1208_;
  assign new_n1210_ = ~controlPi_17_2 & new_n1209_;
  assign new_n1211_ = ~controlPi_17_1 & ~n428_ntk1;
  assign new_n1212_ = controlPi_17_1 & ~n435_ntk1;
  assign new_n1213_ = ~new_n1211_ & ~new_n1212_;
  assign new_n1214_ = controlPi_17_2 & new_n1213_;
  assign new_n1215_ = ~new_n1210_ & ~new_n1214_;
  assign new_n1216_ = controlPi_17_3 & new_n1215_;
  assign new_n1217_ = ~new_n1206_ & ~new_n1216_;
  assign new_n1218_ = controlPi_17_4 & ~new_n1217_;
  assign new_n1219_ = ~controlPi_17_1 & ~n2_ntk1;
  assign new_n1220_ = controlPi_17_1 & ~n13_ntk1;
  assign new_n1221_ = ~new_n1219_ & ~new_n1220_;
  assign new_n1222_ = ~controlPi_17_2 & new_n1221_;
  assign new_n1223_ = ~controlPi_17_1 & ~n46_ntk1;
  assign new_n1224_ = controlPi_17_1 & ~n75_ntk1;
  assign new_n1225_ = ~new_n1223_ & ~new_n1224_;
  assign new_n1226_ = controlPi_17_2 & new_n1225_;
  assign new_n1227_ = ~new_n1222_ & ~new_n1226_;
  assign new_n1228_ = ~controlPi_17_3 & new_n1227_;
  assign new_n1229_ = ~controlPi_17_1 & ~n96_ntk1;
  assign new_n1230_ = controlPi_17_1 & ~n131_ntk1;
  assign new_n1231_ = ~new_n1229_ & ~new_n1230_;
  assign new_n1232_ = ~controlPi_17_2 & new_n1231_;
  assign new_n1233_ = ~controlPi_17_1 & ~n159_ntk1;
  assign new_n1234_ = controlPi_17_1 & ~n177_ntk1;
  assign new_n1235_ = ~new_n1233_ & ~new_n1234_;
  assign new_n1236_ = controlPi_17_2 & new_n1235_;
  assign new_n1237_ = ~new_n1232_ & ~new_n1236_;
  assign new_n1238_ = controlPi_17_3 & new_n1237_;
  assign new_n1239_ = ~new_n1228_ & ~new_n1238_;
  assign new_n1240_ = ~controlPi_17_4 & ~new_n1239_;
  assign new_n1241_ = ~new_n1218_ & ~new_n1240_;
  assign new_n1242_ = ~controlPi_17_5 & ~new_n1241_;
  assign new_n1243_ = controlPi_17_1 & n659_ntk1;
  assign new_n1244_ = ~controlPi_17_1 & n616_ntk1;
  assign new_n1245_ = ~new_n1243_ & ~new_n1244_;
  assign new_n1246_ = ~controlPi_17_2 & new_n1245_;
  assign new_n1247_ = controlPi_17_1 & n673_ntk1;
  assign new_n1248_ = ~controlPi_17_1 & n664_ntk1;
  assign new_n1249_ = ~new_n1247_ & ~new_n1248_;
  assign new_n1250_ = controlPi_17_2 & new_n1249_;
  assign new_n1251_ = ~new_n1246_ & ~new_n1250_;
  assign new_n1252_ = controlPi_17_4 & ~new_n1251_;
  assign new_n1253_ = controlPi_17_1 & n457_ntk1;
  assign new_n1254_ = ~controlPi_17_1 & n454_ntk1;
  assign new_n1255_ = ~new_n1253_ & ~new_n1254_;
  assign new_n1256_ = ~controlPi_17_2 & new_n1255_;
  assign new_n1257_ = controlPi_17_1 & n507_ntk1;
  assign new_n1258_ = ~controlPi_17_1 & n468_ntk1;
  assign new_n1259_ = ~new_n1257_ & ~new_n1258_;
  assign new_n1260_ = controlPi_17_2 & new_n1259_;
  assign new_n1261_ = ~new_n1256_ & ~new_n1260_;
  assign new_n1262_ = ~controlPi_17_4 & ~new_n1261_;
  assign new_n1263_ = ~new_n1252_ & ~new_n1262_;
  assign new_n1264_ = ~controlPi_17_3 & ~new_n1263_;
  assign new_n1265_ = controlPi_17_1 & n600_ntk1;
  assign new_n1266_ = ~controlPi_17_1 & n582_ntk1;
  assign new_n1267_ = ~new_n1265_ & ~new_n1266_;
  assign new_n1268_ = controlPi_17_2 & new_n1267_;
  assign new_n1269_ = controlPi_17_1 & n525_ntk1;
  assign new_n1270_ = ~controlPi_17_1 & n511_ntk1;
  assign new_n1271_ = ~new_n1269_ & ~new_n1270_;
  assign new_n1272_ = ~controlPi_17_2 & new_n1271_;
  assign new_n1273_ = ~new_n1268_ & ~new_n1272_;
  assign new_n1274_ = controlPi_17_3 & ~new_n1273_;
  assign new_n1275_ = ~controlPi_17_4 & new_n1274_;
  assign new_n1276_ = ~new_n1264_ & ~new_n1275_;
  assign new_n1277_ = controlPi_17_5 & ~new_n1276_;
  assign new_n1278_ = ~new_n1242_ & ~new_n1277_;
  assign new_n1279_ = controlPi_17_0 & ~new_n1278_;
  assign new_n1280_ = ~controlPi_17_0 & new_n1278_;
  assign new_n1281_ = ~new_n1279_ & ~new_n1280_;
  assign new_n1282_ = ~controlPi_37_1 & ~n199_ntk1;
  assign new_n1283_ = controlPi_37_1 & ~n211_ntk1;
  assign new_n1284_ = ~new_n1282_ & ~new_n1283_;
  assign new_n1285_ = ~controlPi_37_2 & new_n1284_;
  assign new_n1286_ = ~controlPi_37_1 & ~n216_ntk1;
  assign new_n1287_ = controlPi_37_1 & ~n280_ntk1;
  assign new_n1288_ = ~new_n1286_ & ~new_n1287_;
  assign new_n1289_ = controlPi_37_2 & new_n1288_;
  assign new_n1290_ = ~new_n1285_ & ~new_n1289_;
  assign new_n1291_ = ~controlPi_37_3 & new_n1290_;
  assign new_n1292_ = ~controlPi_37_1 & ~n287_ntk1;
  assign new_n1293_ = controlPi_37_1 & ~n409_ntk1;
  assign new_n1294_ = ~new_n1292_ & ~new_n1293_;
  assign new_n1295_ = ~controlPi_37_2 & new_n1294_;
  assign new_n1296_ = ~controlPi_37_1 & ~n428_ntk1;
  assign new_n1297_ = controlPi_37_1 & ~n435_ntk1;
  assign new_n1298_ = ~new_n1296_ & ~new_n1297_;
  assign new_n1299_ = controlPi_37_2 & new_n1298_;
  assign new_n1300_ = ~new_n1295_ & ~new_n1299_;
  assign new_n1301_ = controlPi_37_3 & new_n1300_;
  assign new_n1302_ = ~new_n1291_ & ~new_n1301_;
  assign new_n1303_ = controlPi_37_4 & ~new_n1302_;
  assign new_n1304_ = ~controlPi_37_1 & ~n2_ntk1;
  assign new_n1305_ = controlPi_37_1 & ~n13_ntk1;
  assign new_n1306_ = ~new_n1304_ & ~new_n1305_;
  assign new_n1307_ = ~controlPi_37_2 & new_n1306_;
  assign new_n1308_ = ~controlPi_37_1 & ~n46_ntk1;
  assign new_n1309_ = controlPi_37_1 & ~n75_ntk1;
  assign new_n1310_ = ~new_n1308_ & ~new_n1309_;
  assign new_n1311_ = controlPi_37_2 & new_n1310_;
  assign new_n1312_ = ~new_n1307_ & ~new_n1311_;
  assign new_n1313_ = ~controlPi_37_3 & new_n1312_;
  assign new_n1314_ = ~controlPi_37_1 & ~n96_ntk1;
  assign new_n1315_ = controlPi_37_1 & ~n131_ntk1;
  assign new_n1316_ = ~new_n1314_ & ~new_n1315_;
  assign new_n1317_ = ~controlPi_37_2 & new_n1316_;
  assign new_n1318_ = ~controlPi_37_1 & ~n159_ntk1;
  assign new_n1319_ = controlPi_37_1 & ~n177_ntk1;
  assign new_n1320_ = ~new_n1318_ & ~new_n1319_;
  assign new_n1321_ = controlPi_37_2 & new_n1320_;
  assign new_n1322_ = ~new_n1317_ & ~new_n1321_;
  assign new_n1323_ = controlPi_37_3 & new_n1322_;
  assign new_n1324_ = ~new_n1313_ & ~new_n1323_;
  assign new_n1325_ = ~controlPi_37_4 & ~new_n1324_;
  assign new_n1326_ = ~new_n1303_ & ~new_n1325_;
  assign new_n1327_ = ~controlPi_37_5 & ~new_n1326_;
  assign new_n1328_ = controlPi_37_1 & n659_ntk1;
  assign new_n1329_ = ~controlPi_37_1 & n616_ntk1;
  assign new_n1330_ = ~new_n1328_ & ~new_n1329_;
  assign new_n1331_ = ~controlPi_37_2 & new_n1330_;
  assign new_n1332_ = controlPi_37_1 & n673_ntk1;
  assign new_n1333_ = ~controlPi_37_1 & n664_ntk1;
  assign new_n1334_ = ~new_n1332_ & ~new_n1333_;
  assign new_n1335_ = controlPi_37_2 & new_n1334_;
  assign new_n1336_ = ~new_n1331_ & ~new_n1335_;
  assign new_n1337_ = controlPi_37_4 & ~new_n1336_;
  assign new_n1338_ = controlPi_37_1 & n457_ntk1;
  assign new_n1339_ = ~controlPi_37_1 & n454_ntk1;
  assign new_n1340_ = ~new_n1338_ & ~new_n1339_;
  assign new_n1341_ = ~controlPi_37_2 & new_n1340_;
  assign new_n1342_ = controlPi_37_1 & n507_ntk1;
  assign new_n1343_ = ~controlPi_37_1 & n468_ntk1;
  assign new_n1344_ = ~new_n1342_ & ~new_n1343_;
  assign new_n1345_ = controlPi_37_2 & new_n1344_;
  assign new_n1346_ = ~new_n1341_ & ~new_n1345_;
  assign new_n1347_ = ~controlPi_37_4 & ~new_n1346_;
  assign new_n1348_ = ~new_n1337_ & ~new_n1347_;
  assign new_n1349_ = ~controlPi_37_3 & ~new_n1348_;
  assign new_n1350_ = controlPi_37_1 & n600_ntk1;
  assign new_n1351_ = ~controlPi_37_1 & n582_ntk1;
  assign new_n1352_ = ~new_n1350_ & ~new_n1351_;
  assign new_n1353_ = controlPi_37_2 & new_n1352_;
  assign new_n1354_ = controlPi_37_1 & n525_ntk1;
  assign new_n1355_ = ~controlPi_37_1 & n511_ntk1;
  assign new_n1356_ = ~new_n1354_ & ~new_n1355_;
  assign new_n1357_ = ~controlPi_37_2 & new_n1356_;
  assign new_n1358_ = ~new_n1353_ & ~new_n1357_;
  assign new_n1359_ = controlPi_37_3 & ~new_n1358_;
  assign new_n1360_ = ~controlPi_37_4 & new_n1359_;
  assign new_n1361_ = ~new_n1349_ & ~new_n1360_;
  assign new_n1362_ = controlPi_37_5 & ~new_n1361_;
  assign new_n1363_ = ~new_n1327_ & ~new_n1362_;
  assign new_n1364_ = controlPi_37_0 & ~new_n1363_;
  assign new_n1365_ = ~controlPi_37_0 & new_n1363_;
  assign new_n1366_ = ~new_n1364_ & ~new_n1365_;
  assign new_n1367_ = ~new_n1281_ & ~new_n1366_;
  assign new_n1368_ = new_n1110_ & new_n1195_;
  assign new_n1369_ = new_n1367_ & ~new_n1368_;
  assign new_n1370_ = ~new_n1196_ & ~new_n1369_;
  assign new_n1371_ = ~controlPi_64_1 & ~n199_ntk1;
  assign new_n1372_ = controlPi_64_1 & ~n211_ntk1;
  assign new_n1373_ = ~new_n1371_ & ~new_n1372_;
  assign new_n1374_ = ~controlPi_64_2 & new_n1373_;
  assign new_n1375_ = ~controlPi_64_1 & ~n216_ntk1;
  assign new_n1376_ = controlPi_64_1 & ~n280_ntk1;
  assign new_n1377_ = ~new_n1375_ & ~new_n1376_;
  assign new_n1378_ = controlPi_64_2 & new_n1377_;
  assign new_n1379_ = ~new_n1374_ & ~new_n1378_;
  assign new_n1380_ = ~controlPi_64_3 & new_n1379_;
  assign new_n1381_ = ~controlPi_64_1 & ~n287_ntk1;
  assign new_n1382_ = controlPi_64_1 & ~n409_ntk1;
  assign new_n1383_ = ~new_n1381_ & ~new_n1382_;
  assign new_n1384_ = ~controlPi_64_2 & new_n1383_;
  assign new_n1385_ = ~controlPi_64_1 & ~n428_ntk1;
  assign new_n1386_ = controlPi_64_1 & ~n435_ntk1;
  assign new_n1387_ = ~new_n1385_ & ~new_n1386_;
  assign new_n1388_ = controlPi_64_2 & new_n1387_;
  assign new_n1389_ = ~new_n1384_ & ~new_n1388_;
  assign new_n1390_ = controlPi_64_3 & new_n1389_;
  assign new_n1391_ = ~new_n1380_ & ~new_n1390_;
  assign new_n1392_ = controlPi_64_4 & ~new_n1391_;
  assign new_n1393_ = ~controlPi_64_1 & ~n2_ntk1;
  assign new_n1394_ = controlPi_64_1 & ~n13_ntk1;
  assign new_n1395_ = ~new_n1393_ & ~new_n1394_;
  assign new_n1396_ = ~controlPi_64_2 & new_n1395_;
  assign new_n1397_ = ~controlPi_64_1 & ~n46_ntk1;
  assign new_n1398_ = controlPi_64_1 & ~n75_ntk1;
  assign new_n1399_ = ~new_n1397_ & ~new_n1398_;
  assign new_n1400_ = controlPi_64_2 & new_n1399_;
  assign new_n1401_ = ~new_n1396_ & ~new_n1400_;
  assign new_n1402_ = ~controlPi_64_3 & new_n1401_;
  assign new_n1403_ = ~controlPi_64_1 & ~n96_ntk1;
  assign new_n1404_ = controlPi_64_1 & ~n131_ntk1;
  assign new_n1405_ = ~new_n1403_ & ~new_n1404_;
  assign new_n1406_ = ~controlPi_64_2 & new_n1405_;
  assign new_n1407_ = ~controlPi_64_1 & ~n159_ntk1;
  assign new_n1408_ = controlPi_64_1 & ~n177_ntk1;
  assign new_n1409_ = ~new_n1407_ & ~new_n1408_;
  assign new_n1410_ = controlPi_64_2 & new_n1409_;
  assign new_n1411_ = ~new_n1406_ & ~new_n1410_;
  assign new_n1412_ = controlPi_64_3 & new_n1411_;
  assign new_n1413_ = ~new_n1402_ & ~new_n1412_;
  assign new_n1414_ = ~controlPi_64_4 & ~new_n1413_;
  assign new_n1415_ = ~new_n1392_ & ~new_n1414_;
  assign new_n1416_ = ~controlPi_64_5 & ~new_n1415_;
  assign new_n1417_ = controlPi_64_1 & n659_ntk1;
  assign new_n1418_ = ~controlPi_64_1 & n616_ntk1;
  assign new_n1419_ = ~new_n1417_ & ~new_n1418_;
  assign new_n1420_ = ~controlPi_64_2 & new_n1419_;
  assign new_n1421_ = controlPi_64_1 & n673_ntk1;
  assign new_n1422_ = ~controlPi_64_1 & n664_ntk1;
  assign new_n1423_ = ~new_n1421_ & ~new_n1422_;
  assign new_n1424_ = controlPi_64_2 & new_n1423_;
  assign new_n1425_ = ~new_n1420_ & ~new_n1424_;
  assign new_n1426_ = controlPi_64_4 & ~new_n1425_;
  assign new_n1427_ = controlPi_64_1 & n457_ntk1;
  assign new_n1428_ = ~controlPi_64_1 & n454_ntk1;
  assign new_n1429_ = ~new_n1427_ & ~new_n1428_;
  assign new_n1430_ = ~controlPi_64_2 & new_n1429_;
  assign new_n1431_ = controlPi_64_1 & n507_ntk1;
  assign new_n1432_ = ~controlPi_64_1 & n468_ntk1;
  assign new_n1433_ = ~new_n1431_ & ~new_n1432_;
  assign new_n1434_ = controlPi_64_2 & new_n1433_;
  assign new_n1435_ = ~new_n1430_ & ~new_n1434_;
  assign new_n1436_ = ~controlPi_64_4 & ~new_n1435_;
  assign new_n1437_ = ~new_n1426_ & ~new_n1436_;
  assign new_n1438_ = ~controlPi_64_3 & ~new_n1437_;
  assign new_n1439_ = controlPi_64_1 & n600_ntk1;
  assign new_n1440_ = ~controlPi_64_1 & n582_ntk1;
  assign new_n1441_ = ~new_n1439_ & ~new_n1440_;
  assign new_n1442_ = controlPi_64_2 & new_n1441_;
  assign new_n1443_ = controlPi_64_1 & n525_ntk1;
  assign new_n1444_ = ~controlPi_64_1 & n511_ntk1;
  assign new_n1445_ = ~new_n1443_ & ~new_n1444_;
  assign new_n1446_ = ~controlPi_64_2 & new_n1445_;
  assign new_n1447_ = ~new_n1442_ & ~new_n1446_;
  assign new_n1448_ = controlPi_64_3 & ~new_n1447_;
  assign new_n1449_ = ~controlPi_64_4 & new_n1448_;
  assign new_n1450_ = ~new_n1438_ & ~new_n1449_;
  assign new_n1451_ = controlPi_64_5 & ~new_n1450_;
  assign new_n1452_ = ~new_n1416_ & ~new_n1451_;
  assign new_n1453_ = controlPi_64_0 & ~new_n1452_;
  assign new_n1454_ = ~controlPi_64_0 & new_n1452_;
  assign new_n1455_ = ~new_n1453_ & ~new_n1454_;
  assign new_n1456_ = ~controlPi_71_1 & ~n199_ntk1;
  assign new_n1457_ = controlPi_71_1 & ~n211_ntk1;
  assign new_n1458_ = ~new_n1456_ & ~new_n1457_;
  assign new_n1459_ = ~controlPi_71_2 & new_n1458_;
  assign new_n1460_ = ~controlPi_71_1 & ~n216_ntk1;
  assign new_n1461_ = controlPi_71_1 & ~n280_ntk1;
  assign new_n1462_ = ~new_n1460_ & ~new_n1461_;
  assign new_n1463_ = controlPi_71_2 & new_n1462_;
  assign new_n1464_ = ~new_n1459_ & ~new_n1463_;
  assign new_n1465_ = ~controlPi_71_3 & new_n1464_;
  assign new_n1466_ = ~controlPi_71_1 & ~n287_ntk1;
  assign new_n1467_ = controlPi_71_1 & ~n409_ntk1;
  assign new_n1468_ = ~new_n1466_ & ~new_n1467_;
  assign new_n1469_ = ~controlPi_71_2 & new_n1468_;
  assign new_n1470_ = ~controlPi_71_1 & ~n428_ntk1;
  assign new_n1471_ = controlPi_71_1 & ~n435_ntk1;
  assign new_n1472_ = ~new_n1470_ & ~new_n1471_;
  assign new_n1473_ = controlPi_71_2 & new_n1472_;
  assign new_n1474_ = ~new_n1469_ & ~new_n1473_;
  assign new_n1475_ = controlPi_71_3 & new_n1474_;
  assign new_n1476_ = ~new_n1465_ & ~new_n1475_;
  assign new_n1477_ = controlPi_71_4 & ~new_n1476_;
  assign new_n1478_ = ~controlPi_71_1 & ~n2_ntk1;
  assign new_n1479_ = controlPi_71_1 & ~n13_ntk1;
  assign new_n1480_ = ~new_n1478_ & ~new_n1479_;
  assign new_n1481_ = ~controlPi_71_2 & new_n1480_;
  assign new_n1482_ = ~controlPi_71_1 & ~n46_ntk1;
  assign new_n1483_ = controlPi_71_1 & ~n75_ntk1;
  assign new_n1484_ = ~new_n1482_ & ~new_n1483_;
  assign new_n1485_ = controlPi_71_2 & new_n1484_;
  assign new_n1486_ = ~new_n1481_ & ~new_n1485_;
  assign new_n1487_ = ~controlPi_71_3 & new_n1486_;
  assign new_n1488_ = ~controlPi_71_1 & ~n96_ntk1;
  assign new_n1489_ = controlPi_71_1 & ~n131_ntk1;
  assign new_n1490_ = ~new_n1488_ & ~new_n1489_;
  assign new_n1491_ = ~controlPi_71_2 & new_n1490_;
  assign new_n1492_ = ~controlPi_71_1 & ~n159_ntk1;
  assign new_n1493_ = controlPi_71_1 & ~n177_ntk1;
  assign new_n1494_ = ~new_n1492_ & ~new_n1493_;
  assign new_n1495_ = controlPi_71_2 & new_n1494_;
  assign new_n1496_ = ~new_n1491_ & ~new_n1495_;
  assign new_n1497_ = controlPi_71_3 & new_n1496_;
  assign new_n1498_ = ~new_n1487_ & ~new_n1497_;
  assign new_n1499_ = ~controlPi_71_4 & ~new_n1498_;
  assign new_n1500_ = ~new_n1477_ & ~new_n1499_;
  assign new_n1501_ = ~controlPi_71_5 & ~new_n1500_;
  assign new_n1502_ = controlPi_71_1 & n659_ntk1;
  assign new_n1503_ = ~controlPi_71_1 & n616_ntk1;
  assign new_n1504_ = ~new_n1502_ & ~new_n1503_;
  assign new_n1505_ = ~controlPi_71_2 & new_n1504_;
  assign new_n1506_ = controlPi_71_1 & n673_ntk1;
  assign new_n1507_ = ~controlPi_71_1 & n664_ntk1;
  assign new_n1508_ = ~new_n1506_ & ~new_n1507_;
  assign new_n1509_ = controlPi_71_2 & new_n1508_;
  assign new_n1510_ = ~new_n1505_ & ~new_n1509_;
  assign new_n1511_ = controlPi_71_4 & ~new_n1510_;
  assign new_n1512_ = controlPi_71_1 & n457_ntk1;
  assign new_n1513_ = ~controlPi_71_1 & n454_ntk1;
  assign new_n1514_ = ~new_n1512_ & ~new_n1513_;
  assign new_n1515_ = ~controlPi_71_2 & new_n1514_;
  assign new_n1516_ = controlPi_71_1 & n507_ntk1;
  assign new_n1517_ = ~controlPi_71_1 & n468_ntk1;
  assign new_n1518_ = ~new_n1516_ & ~new_n1517_;
  assign new_n1519_ = controlPi_71_2 & new_n1518_;
  assign new_n1520_ = ~new_n1515_ & ~new_n1519_;
  assign new_n1521_ = ~controlPi_71_4 & ~new_n1520_;
  assign new_n1522_ = ~new_n1511_ & ~new_n1521_;
  assign new_n1523_ = ~controlPi_71_3 & ~new_n1522_;
  assign new_n1524_ = controlPi_71_1 & n600_ntk1;
  assign new_n1525_ = ~controlPi_71_1 & n582_ntk1;
  assign new_n1526_ = ~new_n1524_ & ~new_n1525_;
  assign new_n1527_ = controlPi_71_2 & new_n1526_;
  assign new_n1528_ = controlPi_71_1 & n525_ntk1;
  assign new_n1529_ = ~controlPi_71_1 & n511_ntk1;
  assign new_n1530_ = ~new_n1528_ & ~new_n1529_;
  assign new_n1531_ = ~controlPi_71_2 & new_n1530_;
  assign new_n1532_ = ~new_n1527_ & ~new_n1531_;
  assign new_n1533_ = controlPi_71_3 & ~new_n1532_;
  assign new_n1534_ = ~controlPi_71_4 & new_n1533_;
  assign new_n1535_ = ~new_n1523_ & ~new_n1534_;
  assign new_n1536_ = controlPi_71_5 & ~new_n1535_;
  assign new_n1537_ = ~new_n1501_ & ~new_n1536_;
  assign new_n1538_ = controlPi_71_0 & ~new_n1537_;
  assign new_n1539_ = ~controlPi_71_0 & new_n1537_;
  assign new_n1540_ = ~new_n1538_ & ~new_n1539_;
  assign new_n1541_ = ~new_n1455_ & ~new_n1540_;
  assign new_n1542_ = new_n1455_ & new_n1540_;
  assign new_n1543_ = ~new_n1541_ & ~new_n1542_;
  assign new_n1544_ = new_n1370_ & ~new_n1543_;
  assign new_n1545_ = ~new_n1370_ & new_n1543_;
  assign new_n1546_ = ~new_n939_ & ~new_n1545_;
  assign new_n1547_ = ~new_n1544_ & new_n1546_;
  assign new_n1548_ = ~new_n1025_ & ~new_n1547_;
  assign new_n1549_ = ~controlPi_44_1 & ~n349_ntk1;
  assign new_n1550_ = controlPi_44_1 & ~n368_ntk1;
  assign new_n1551_ = ~new_n1549_ & ~new_n1550_;
  assign new_n1552_ = controlPi_44_3 & ~new_n1551_;
  assign new_n1553_ = ~controlPi_44_1 & ~n85_ntk1;
  assign new_n1554_ = controlPi_44_1 & ~n93_ntk1;
  assign new_n1555_ = ~new_n1553_ & ~new_n1554_;
  assign new_n1556_ = ~controlPi_44_3 & ~new_n1555_;
  assign new_n1557_ = ~new_n1552_ & ~new_n1556_;
  assign new_n1558_ = ~controlPi_44_2 & ~new_n1557_;
  assign new_n1559_ = ~controlPi_44_1 & ~n206_ntk1;
  assign new_n1560_ = controlPi_44_1 & ~n266_ntk1;
  assign new_n1561_ = ~new_n1559_ & ~new_n1560_;
  assign new_n1562_ = controlPi_44_2 & ~new_n1561_;
  assign new_n1563_ = ~controlPi_44_3 & new_n1562_;
  assign new_n1564_ = ~new_n1558_ & ~new_n1563_;
  assign new_n1565_ = controlPi_44_0 & ~new_n1564_;
  assign new_n1566_ = ~controlPi_44_0 & new_n1564_;
  assign new_n1567_ = ~new_n1565_ & ~new_n1566_;
  assign new_n1568_ = ~controlPi_45_1 & ~n349_ntk1;
  assign new_n1569_ = controlPi_45_1 & ~n368_ntk1;
  assign new_n1570_ = ~new_n1568_ & ~new_n1569_;
  assign new_n1571_ = controlPi_45_3 & ~new_n1570_;
  assign new_n1572_ = ~controlPi_45_1 & ~n85_ntk1;
  assign new_n1573_ = controlPi_45_1 & ~n93_ntk1;
  assign new_n1574_ = ~new_n1572_ & ~new_n1573_;
  assign new_n1575_ = ~controlPi_45_3 & ~new_n1574_;
  assign new_n1576_ = ~new_n1571_ & ~new_n1575_;
  assign new_n1577_ = ~controlPi_45_2 & ~new_n1576_;
  assign new_n1578_ = ~controlPi_45_1 & ~n206_ntk1;
  assign new_n1579_ = controlPi_45_1 & ~n266_ntk1;
  assign new_n1580_ = ~new_n1578_ & ~new_n1579_;
  assign new_n1581_ = controlPi_45_2 & ~new_n1580_;
  assign new_n1582_ = ~controlPi_45_3 & new_n1581_;
  assign new_n1583_ = ~new_n1577_ & ~new_n1582_;
  assign new_n1584_ = controlPi_45_0 & ~new_n1583_;
  assign new_n1585_ = ~controlPi_45_0 & new_n1583_;
  assign new_n1586_ = ~new_n1584_ & ~new_n1585_;
  assign new_n1587_ = ~controlPi_60_1 & ~n349_ntk1;
  assign new_n1588_ = controlPi_60_1 & ~n368_ntk1;
  assign new_n1589_ = ~new_n1587_ & ~new_n1588_;
  assign new_n1590_ = controlPi_60_3 & ~new_n1589_;
  assign new_n1591_ = ~controlPi_60_1 & ~n85_ntk1;
  assign new_n1592_ = controlPi_60_1 & ~n93_ntk1;
  assign new_n1593_ = ~new_n1591_ & ~new_n1592_;
  assign new_n1594_ = ~controlPi_60_3 & ~new_n1593_;
  assign new_n1595_ = ~new_n1590_ & ~new_n1594_;
  assign new_n1596_ = ~controlPi_60_2 & ~new_n1595_;
  assign new_n1597_ = ~controlPi_60_1 & ~n206_ntk1;
  assign new_n1598_ = controlPi_60_1 & ~n266_ntk1;
  assign new_n1599_ = ~new_n1597_ & ~new_n1598_;
  assign new_n1600_ = controlPi_60_2 & ~new_n1599_;
  assign new_n1601_ = ~controlPi_60_3 & new_n1600_;
  assign new_n1602_ = ~new_n1596_ & ~new_n1601_;
  assign new_n1603_ = controlPi_60_0 & ~new_n1602_;
  assign new_n1604_ = ~controlPi_60_0 & new_n1602_;
  assign new_n1605_ = ~new_n1603_ & ~new_n1604_;
  assign new_n1606_ = ~controlPi_32_1 & ~n199_ntk1;
  assign new_n1607_ = controlPi_32_1 & ~n211_ntk1;
  assign new_n1608_ = ~new_n1606_ & ~new_n1607_;
  assign new_n1609_ = ~controlPi_32_2 & new_n1608_;
  assign new_n1610_ = ~controlPi_32_1 & ~n216_ntk1;
  assign new_n1611_ = controlPi_32_1 & ~n280_ntk1;
  assign new_n1612_ = ~new_n1610_ & ~new_n1611_;
  assign new_n1613_ = controlPi_32_2 & new_n1612_;
  assign new_n1614_ = ~new_n1609_ & ~new_n1613_;
  assign new_n1615_ = ~controlPi_32_3 & new_n1614_;
  assign new_n1616_ = ~controlPi_32_1 & ~n287_ntk1;
  assign new_n1617_ = controlPi_32_1 & ~n409_ntk1;
  assign new_n1618_ = ~new_n1616_ & ~new_n1617_;
  assign new_n1619_ = ~controlPi_32_2 & new_n1618_;
  assign new_n1620_ = ~controlPi_32_1 & ~n428_ntk1;
  assign new_n1621_ = controlPi_32_1 & ~n435_ntk1;
  assign new_n1622_ = ~new_n1620_ & ~new_n1621_;
  assign new_n1623_ = controlPi_32_2 & new_n1622_;
  assign new_n1624_ = ~new_n1619_ & ~new_n1623_;
  assign new_n1625_ = controlPi_32_3 & new_n1624_;
  assign new_n1626_ = ~new_n1615_ & ~new_n1625_;
  assign new_n1627_ = controlPi_32_4 & ~new_n1626_;
  assign new_n1628_ = ~controlPi_32_1 & ~n2_ntk1;
  assign new_n1629_ = controlPi_32_1 & ~n13_ntk1;
  assign new_n1630_ = ~new_n1628_ & ~new_n1629_;
  assign new_n1631_ = ~controlPi_32_2 & new_n1630_;
  assign new_n1632_ = ~controlPi_32_1 & ~n46_ntk1;
  assign new_n1633_ = controlPi_32_1 & ~n75_ntk1;
  assign new_n1634_ = ~new_n1632_ & ~new_n1633_;
  assign new_n1635_ = controlPi_32_2 & new_n1634_;
  assign new_n1636_ = ~new_n1631_ & ~new_n1635_;
  assign new_n1637_ = ~controlPi_32_3 & new_n1636_;
  assign new_n1638_ = ~controlPi_32_1 & ~n96_ntk1;
  assign new_n1639_ = controlPi_32_1 & ~n131_ntk1;
  assign new_n1640_ = ~new_n1638_ & ~new_n1639_;
  assign new_n1641_ = ~controlPi_32_2 & new_n1640_;
  assign new_n1642_ = ~controlPi_32_1 & ~n159_ntk1;
  assign new_n1643_ = controlPi_32_1 & ~n177_ntk1;
  assign new_n1644_ = ~new_n1642_ & ~new_n1643_;
  assign new_n1645_ = controlPi_32_2 & new_n1644_;
  assign new_n1646_ = ~new_n1641_ & ~new_n1645_;
  assign new_n1647_ = controlPi_32_3 & new_n1646_;
  assign new_n1648_ = ~new_n1637_ & ~new_n1647_;
  assign new_n1649_ = ~controlPi_32_4 & ~new_n1648_;
  assign new_n1650_ = ~new_n1627_ & ~new_n1649_;
  assign new_n1651_ = ~controlPi_32_5 & ~new_n1650_;
  assign new_n1652_ = controlPi_32_1 & n659_ntk1;
  assign new_n1653_ = ~controlPi_32_1 & n616_ntk1;
  assign new_n1654_ = ~new_n1652_ & ~new_n1653_;
  assign new_n1655_ = ~controlPi_32_2 & new_n1654_;
  assign new_n1656_ = controlPi_32_1 & n673_ntk1;
  assign new_n1657_ = ~controlPi_32_1 & n664_ntk1;
  assign new_n1658_ = ~new_n1656_ & ~new_n1657_;
  assign new_n1659_ = controlPi_32_2 & new_n1658_;
  assign new_n1660_ = ~new_n1655_ & ~new_n1659_;
  assign new_n1661_ = controlPi_32_4 & ~new_n1660_;
  assign new_n1662_ = controlPi_32_1 & n457_ntk1;
  assign new_n1663_ = ~controlPi_32_1 & n454_ntk1;
  assign new_n1664_ = ~new_n1662_ & ~new_n1663_;
  assign new_n1665_ = ~controlPi_32_2 & new_n1664_;
  assign new_n1666_ = controlPi_32_1 & n507_ntk1;
  assign new_n1667_ = ~controlPi_32_1 & n468_ntk1;
  assign new_n1668_ = ~new_n1666_ & ~new_n1667_;
  assign new_n1669_ = controlPi_32_2 & new_n1668_;
  assign new_n1670_ = ~new_n1665_ & ~new_n1669_;
  assign new_n1671_ = ~controlPi_32_4 & ~new_n1670_;
  assign new_n1672_ = ~new_n1661_ & ~new_n1671_;
  assign new_n1673_ = ~controlPi_32_3 & ~new_n1672_;
  assign new_n1674_ = controlPi_32_1 & n600_ntk1;
  assign new_n1675_ = ~controlPi_32_1 & n582_ntk1;
  assign new_n1676_ = ~new_n1674_ & ~new_n1675_;
  assign new_n1677_ = controlPi_32_2 & new_n1676_;
  assign new_n1678_ = controlPi_32_1 & n525_ntk1;
  assign new_n1679_ = ~controlPi_32_1 & n511_ntk1;
  assign new_n1680_ = ~new_n1678_ & ~new_n1679_;
  assign new_n1681_ = ~controlPi_32_2 & new_n1680_;
  assign new_n1682_ = ~new_n1677_ & ~new_n1681_;
  assign new_n1683_ = controlPi_32_3 & ~new_n1682_;
  assign new_n1684_ = ~controlPi_32_4 & new_n1683_;
  assign new_n1685_ = ~new_n1673_ & ~new_n1684_;
  assign new_n1686_ = controlPi_32_5 & ~new_n1685_;
  assign new_n1687_ = ~new_n1651_ & ~new_n1686_;
  assign new_n1688_ = controlPi_32_0 & ~new_n1687_;
  assign new_n1689_ = ~controlPi_32_0 & new_n1687_;
  assign new_n1690_ = ~new_n1688_ & ~new_n1689_;
  assign new_n1691_ = ~controlPi_49_1 & ~n199_ntk1;
  assign new_n1692_ = controlPi_49_1 & ~n211_ntk1;
  assign new_n1693_ = ~new_n1691_ & ~new_n1692_;
  assign new_n1694_ = ~controlPi_49_2 & new_n1693_;
  assign new_n1695_ = ~controlPi_49_1 & ~n216_ntk1;
  assign new_n1696_ = controlPi_49_1 & ~n280_ntk1;
  assign new_n1697_ = ~new_n1695_ & ~new_n1696_;
  assign new_n1698_ = controlPi_49_2 & new_n1697_;
  assign new_n1699_ = ~new_n1694_ & ~new_n1698_;
  assign new_n1700_ = ~controlPi_49_3 & new_n1699_;
  assign new_n1701_ = ~controlPi_49_1 & ~n287_ntk1;
  assign new_n1702_ = controlPi_49_1 & ~n409_ntk1;
  assign new_n1703_ = ~new_n1701_ & ~new_n1702_;
  assign new_n1704_ = ~controlPi_49_2 & new_n1703_;
  assign new_n1705_ = ~controlPi_49_1 & ~n428_ntk1;
  assign new_n1706_ = controlPi_49_1 & ~n435_ntk1;
  assign new_n1707_ = ~new_n1705_ & ~new_n1706_;
  assign new_n1708_ = controlPi_49_2 & new_n1707_;
  assign new_n1709_ = ~new_n1704_ & ~new_n1708_;
  assign new_n1710_ = controlPi_49_3 & new_n1709_;
  assign new_n1711_ = ~new_n1700_ & ~new_n1710_;
  assign new_n1712_ = controlPi_49_4 & ~new_n1711_;
  assign new_n1713_ = ~controlPi_49_1 & ~n2_ntk1;
  assign new_n1714_ = controlPi_49_1 & ~n13_ntk1;
  assign new_n1715_ = ~new_n1713_ & ~new_n1714_;
  assign new_n1716_ = ~controlPi_49_2 & new_n1715_;
  assign new_n1717_ = ~controlPi_49_1 & ~n46_ntk1;
  assign new_n1718_ = controlPi_49_1 & ~n75_ntk1;
  assign new_n1719_ = ~new_n1717_ & ~new_n1718_;
  assign new_n1720_ = controlPi_49_2 & new_n1719_;
  assign new_n1721_ = ~new_n1716_ & ~new_n1720_;
  assign new_n1722_ = ~controlPi_49_3 & new_n1721_;
  assign new_n1723_ = ~controlPi_49_1 & ~n96_ntk1;
  assign new_n1724_ = controlPi_49_1 & ~n131_ntk1;
  assign new_n1725_ = ~new_n1723_ & ~new_n1724_;
  assign new_n1726_ = ~controlPi_49_2 & new_n1725_;
  assign new_n1727_ = ~controlPi_49_1 & ~n159_ntk1;
  assign new_n1728_ = controlPi_49_1 & ~n177_ntk1;
  assign new_n1729_ = ~new_n1727_ & ~new_n1728_;
  assign new_n1730_ = controlPi_49_2 & new_n1729_;
  assign new_n1731_ = ~new_n1726_ & ~new_n1730_;
  assign new_n1732_ = controlPi_49_3 & new_n1731_;
  assign new_n1733_ = ~new_n1722_ & ~new_n1732_;
  assign new_n1734_ = ~controlPi_49_4 & ~new_n1733_;
  assign new_n1735_ = ~new_n1712_ & ~new_n1734_;
  assign new_n1736_ = ~controlPi_49_5 & ~new_n1735_;
  assign new_n1737_ = controlPi_49_1 & n659_ntk1;
  assign new_n1738_ = ~controlPi_49_1 & n616_ntk1;
  assign new_n1739_ = ~new_n1737_ & ~new_n1738_;
  assign new_n1740_ = ~controlPi_49_2 & new_n1739_;
  assign new_n1741_ = controlPi_49_1 & n673_ntk1;
  assign new_n1742_ = ~controlPi_49_1 & n664_ntk1;
  assign new_n1743_ = ~new_n1741_ & ~new_n1742_;
  assign new_n1744_ = controlPi_49_2 & new_n1743_;
  assign new_n1745_ = ~new_n1740_ & ~new_n1744_;
  assign new_n1746_ = controlPi_49_4 & ~new_n1745_;
  assign new_n1747_ = controlPi_49_1 & n457_ntk1;
  assign new_n1748_ = ~controlPi_49_1 & n454_ntk1;
  assign new_n1749_ = ~new_n1747_ & ~new_n1748_;
  assign new_n1750_ = ~controlPi_49_2 & new_n1749_;
  assign new_n1751_ = controlPi_49_1 & n507_ntk1;
  assign new_n1752_ = ~controlPi_49_1 & n468_ntk1;
  assign new_n1753_ = ~new_n1751_ & ~new_n1752_;
  assign new_n1754_ = controlPi_49_2 & new_n1753_;
  assign new_n1755_ = ~new_n1750_ & ~new_n1754_;
  assign new_n1756_ = ~controlPi_49_4 & ~new_n1755_;
  assign new_n1757_ = ~new_n1746_ & ~new_n1756_;
  assign new_n1758_ = ~controlPi_49_3 & ~new_n1757_;
  assign new_n1759_ = controlPi_49_1 & n600_ntk1;
  assign new_n1760_ = ~controlPi_49_1 & n582_ntk1;
  assign new_n1761_ = ~new_n1759_ & ~new_n1760_;
  assign new_n1762_ = controlPi_49_2 & new_n1761_;
  assign new_n1763_ = controlPi_49_1 & n525_ntk1;
  assign new_n1764_ = ~controlPi_49_1 & n511_ntk1;
  assign new_n1765_ = ~new_n1763_ & ~new_n1764_;
  assign new_n1766_ = ~controlPi_49_2 & new_n1765_;
  assign new_n1767_ = ~new_n1762_ & ~new_n1766_;
  assign new_n1768_ = controlPi_49_3 & ~new_n1767_;
  assign new_n1769_ = ~controlPi_49_4 & new_n1768_;
  assign new_n1770_ = ~new_n1758_ & ~new_n1769_;
  assign new_n1771_ = controlPi_49_5 & ~new_n1770_;
  assign new_n1772_ = ~new_n1736_ & ~new_n1771_;
  assign new_n1773_ = controlPi_49_0 & ~new_n1772_;
  assign new_n1774_ = ~controlPi_49_0 & new_n1772_;
  assign new_n1775_ = ~new_n1773_ & ~new_n1774_;
  assign new_n1776_ = ~new_n1690_ & ~new_n1775_;
  assign new_n1777_ = ~controlPi_46_1 & ~n199_ntk1;
  assign new_n1778_ = controlPi_46_1 & ~n211_ntk1;
  assign new_n1779_ = ~new_n1777_ & ~new_n1778_;
  assign new_n1780_ = ~controlPi_46_2 & new_n1779_;
  assign new_n1781_ = ~controlPi_46_1 & ~n216_ntk1;
  assign new_n1782_ = controlPi_46_1 & ~n280_ntk1;
  assign new_n1783_ = ~new_n1781_ & ~new_n1782_;
  assign new_n1784_ = controlPi_46_2 & new_n1783_;
  assign new_n1785_ = ~new_n1780_ & ~new_n1784_;
  assign new_n1786_ = ~controlPi_46_3 & new_n1785_;
  assign new_n1787_ = ~controlPi_46_1 & ~n287_ntk1;
  assign new_n1788_ = controlPi_46_1 & ~n409_ntk1;
  assign new_n1789_ = ~new_n1787_ & ~new_n1788_;
  assign new_n1790_ = ~controlPi_46_2 & new_n1789_;
  assign new_n1791_ = ~controlPi_46_1 & ~n428_ntk1;
  assign new_n1792_ = controlPi_46_1 & ~n435_ntk1;
  assign new_n1793_ = ~new_n1791_ & ~new_n1792_;
  assign new_n1794_ = controlPi_46_2 & new_n1793_;
  assign new_n1795_ = ~new_n1790_ & ~new_n1794_;
  assign new_n1796_ = controlPi_46_3 & new_n1795_;
  assign new_n1797_ = ~new_n1786_ & ~new_n1796_;
  assign new_n1798_ = controlPi_46_4 & ~new_n1797_;
  assign new_n1799_ = ~controlPi_46_1 & ~n2_ntk1;
  assign new_n1800_ = controlPi_46_1 & ~n13_ntk1;
  assign new_n1801_ = ~new_n1799_ & ~new_n1800_;
  assign new_n1802_ = ~controlPi_46_2 & new_n1801_;
  assign new_n1803_ = ~controlPi_46_1 & ~n46_ntk1;
  assign new_n1804_ = controlPi_46_1 & ~n75_ntk1;
  assign new_n1805_ = ~new_n1803_ & ~new_n1804_;
  assign new_n1806_ = controlPi_46_2 & new_n1805_;
  assign new_n1807_ = ~new_n1802_ & ~new_n1806_;
  assign new_n1808_ = ~controlPi_46_3 & new_n1807_;
  assign new_n1809_ = ~controlPi_46_1 & ~n96_ntk1;
  assign new_n1810_ = controlPi_46_1 & ~n131_ntk1;
  assign new_n1811_ = ~new_n1809_ & ~new_n1810_;
  assign new_n1812_ = ~controlPi_46_2 & new_n1811_;
  assign new_n1813_ = ~controlPi_46_1 & ~n159_ntk1;
  assign new_n1814_ = controlPi_46_1 & ~n177_ntk1;
  assign new_n1815_ = ~new_n1813_ & ~new_n1814_;
  assign new_n1816_ = controlPi_46_2 & new_n1815_;
  assign new_n1817_ = ~new_n1812_ & ~new_n1816_;
  assign new_n1818_ = controlPi_46_3 & new_n1817_;
  assign new_n1819_ = ~new_n1808_ & ~new_n1818_;
  assign new_n1820_ = ~controlPi_46_4 & ~new_n1819_;
  assign new_n1821_ = ~new_n1798_ & ~new_n1820_;
  assign new_n1822_ = ~controlPi_46_5 & ~new_n1821_;
  assign new_n1823_ = controlPi_46_1 & n659_ntk1;
  assign new_n1824_ = ~controlPi_46_1 & n616_ntk1;
  assign new_n1825_ = ~new_n1823_ & ~new_n1824_;
  assign new_n1826_ = ~controlPi_46_2 & new_n1825_;
  assign new_n1827_ = controlPi_46_1 & n673_ntk1;
  assign new_n1828_ = ~controlPi_46_1 & n664_ntk1;
  assign new_n1829_ = ~new_n1827_ & ~new_n1828_;
  assign new_n1830_ = controlPi_46_2 & new_n1829_;
  assign new_n1831_ = ~new_n1826_ & ~new_n1830_;
  assign new_n1832_ = controlPi_46_4 & ~new_n1831_;
  assign new_n1833_ = controlPi_46_1 & n457_ntk1;
  assign new_n1834_ = ~controlPi_46_1 & n454_ntk1;
  assign new_n1835_ = ~new_n1833_ & ~new_n1834_;
  assign new_n1836_ = ~controlPi_46_2 & new_n1835_;
  assign new_n1837_ = controlPi_46_1 & n507_ntk1;
  assign new_n1838_ = ~controlPi_46_1 & n468_ntk1;
  assign new_n1839_ = ~new_n1837_ & ~new_n1838_;
  assign new_n1840_ = controlPi_46_2 & new_n1839_;
  assign new_n1841_ = ~new_n1836_ & ~new_n1840_;
  assign new_n1842_ = ~controlPi_46_4 & ~new_n1841_;
  assign new_n1843_ = ~new_n1832_ & ~new_n1842_;
  assign new_n1844_ = ~controlPi_46_3 & ~new_n1843_;
  assign new_n1845_ = controlPi_46_1 & n600_ntk1;
  assign new_n1846_ = ~controlPi_46_1 & n582_ntk1;
  assign new_n1847_ = ~new_n1845_ & ~new_n1846_;
  assign new_n1848_ = controlPi_46_2 & new_n1847_;
  assign new_n1849_ = controlPi_46_1 & n525_ntk1;
  assign new_n1850_ = ~controlPi_46_1 & n511_ntk1;
  assign new_n1851_ = ~new_n1849_ & ~new_n1850_;
  assign new_n1852_ = ~controlPi_46_2 & new_n1851_;
  assign new_n1853_ = ~new_n1848_ & ~new_n1852_;
  assign new_n1854_ = controlPi_46_3 & ~new_n1853_;
  assign new_n1855_ = ~controlPi_46_4 & new_n1854_;
  assign new_n1856_ = ~new_n1844_ & ~new_n1855_;
  assign new_n1857_ = controlPi_46_5 & ~new_n1856_;
  assign new_n1858_ = ~new_n1822_ & ~new_n1857_;
  assign new_n1859_ = controlPi_46_0 & ~new_n1858_;
  assign new_n1860_ = ~controlPi_46_0 & new_n1858_;
  assign new_n1861_ = ~new_n1859_ & ~new_n1860_;
  assign new_n1862_ = ~controlPi_67_1 & ~n199_ntk1;
  assign new_n1863_ = controlPi_67_1 & ~n211_ntk1;
  assign new_n1864_ = ~new_n1862_ & ~new_n1863_;
  assign new_n1865_ = ~controlPi_67_2 & new_n1864_;
  assign new_n1866_ = ~controlPi_67_1 & ~n216_ntk1;
  assign new_n1867_ = controlPi_67_1 & ~n280_ntk1;
  assign new_n1868_ = ~new_n1866_ & ~new_n1867_;
  assign new_n1869_ = controlPi_67_2 & new_n1868_;
  assign new_n1870_ = ~new_n1865_ & ~new_n1869_;
  assign new_n1871_ = ~controlPi_67_3 & new_n1870_;
  assign new_n1872_ = ~controlPi_67_1 & ~n287_ntk1;
  assign new_n1873_ = controlPi_67_1 & ~n409_ntk1;
  assign new_n1874_ = ~new_n1872_ & ~new_n1873_;
  assign new_n1875_ = ~controlPi_67_2 & new_n1874_;
  assign new_n1876_ = ~controlPi_67_1 & ~n428_ntk1;
  assign new_n1877_ = controlPi_67_1 & ~n435_ntk1;
  assign new_n1878_ = ~new_n1876_ & ~new_n1877_;
  assign new_n1879_ = controlPi_67_2 & new_n1878_;
  assign new_n1880_ = ~new_n1875_ & ~new_n1879_;
  assign new_n1881_ = controlPi_67_3 & new_n1880_;
  assign new_n1882_ = ~new_n1871_ & ~new_n1881_;
  assign new_n1883_ = controlPi_67_4 & ~new_n1882_;
  assign new_n1884_ = ~controlPi_67_1 & ~n2_ntk1;
  assign new_n1885_ = controlPi_67_1 & ~n13_ntk1;
  assign new_n1886_ = ~new_n1884_ & ~new_n1885_;
  assign new_n1887_ = ~controlPi_67_2 & new_n1886_;
  assign new_n1888_ = ~controlPi_67_1 & ~n46_ntk1;
  assign new_n1889_ = controlPi_67_1 & ~n75_ntk1;
  assign new_n1890_ = ~new_n1888_ & ~new_n1889_;
  assign new_n1891_ = controlPi_67_2 & new_n1890_;
  assign new_n1892_ = ~new_n1887_ & ~new_n1891_;
  assign new_n1893_ = ~controlPi_67_3 & new_n1892_;
  assign new_n1894_ = ~controlPi_67_1 & ~n96_ntk1;
  assign new_n1895_ = controlPi_67_1 & ~n131_ntk1;
  assign new_n1896_ = ~new_n1894_ & ~new_n1895_;
  assign new_n1897_ = ~controlPi_67_2 & new_n1896_;
  assign new_n1898_ = ~controlPi_67_1 & ~n159_ntk1;
  assign new_n1899_ = controlPi_67_1 & ~n177_ntk1;
  assign new_n1900_ = ~new_n1898_ & ~new_n1899_;
  assign new_n1901_ = controlPi_67_2 & new_n1900_;
  assign new_n1902_ = ~new_n1897_ & ~new_n1901_;
  assign new_n1903_ = controlPi_67_3 & new_n1902_;
  assign new_n1904_ = ~new_n1893_ & ~new_n1903_;
  assign new_n1905_ = ~controlPi_67_4 & ~new_n1904_;
  assign new_n1906_ = ~new_n1883_ & ~new_n1905_;
  assign new_n1907_ = ~controlPi_67_5 & ~new_n1906_;
  assign new_n1908_ = controlPi_67_1 & n659_ntk1;
  assign new_n1909_ = ~controlPi_67_1 & n616_ntk1;
  assign new_n1910_ = ~new_n1908_ & ~new_n1909_;
  assign new_n1911_ = ~controlPi_67_2 & new_n1910_;
  assign new_n1912_ = controlPi_67_1 & n673_ntk1;
  assign new_n1913_ = ~controlPi_67_1 & n664_ntk1;
  assign new_n1914_ = ~new_n1912_ & ~new_n1913_;
  assign new_n1915_ = controlPi_67_2 & new_n1914_;
  assign new_n1916_ = ~new_n1911_ & ~new_n1915_;
  assign new_n1917_ = controlPi_67_4 & ~new_n1916_;
  assign new_n1918_ = controlPi_67_1 & n457_ntk1;
  assign new_n1919_ = ~controlPi_67_1 & n454_ntk1;
  assign new_n1920_ = ~new_n1918_ & ~new_n1919_;
  assign new_n1921_ = ~controlPi_67_2 & new_n1920_;
  assign new_n1922_ = controlPi_67_1 & n507_ntk1;
  assign new_n1923_ = ~controlPi_67_1 & n468_ntk1;
  assign new_n1924_ = ~new_n1922_ & ~new_n1923_;
  assign new_n1925_ = controlPi_67_2 & new_n1924_;
  assign new_n1926_ = ~new_n1921_ & ~new_n1925_;
  assign new_n1927_ = ~controlPi_67_4 & ~new_n1926_;
  assign new_n1928_ = ~new_n1917_ & ~new_n1927_;
  assign new_n1929_ = ~controlPi_67_3 & ~new_n1928_;
  assign new_n1930_ = controlPi_67_1 & n600_ntk1;
  assign new_n1931_ = ~controlPi_67_1 & n582_ntk1;
  assign new_n1932_ = ~new_n1930_ & ~new_n1931_;
  assign new_n1933_ = controlPi_67_2 & new_n1932_;
  assign new_n1934_ = controlPi_67_1 & n525_ntk1;
  assign new_n1935_ = ~controlPi_67_1 & n511_ntk1;
  assign new_n1936_ = ~new_n1934_ & ~new_n1935_;
  assign new_n1937_ = ~controlPi_67_2 & new_n1936_;
  assign new_n1938_ = ~new_n1933_ & ~new_n1937_;
  assign new_n1939_ = controlPi_67_3 & ~new_n1938_;
  assign new_n1940_ = ~controlPi_67_4 & new_n1939_;
  assign new_n1941_ = ~new_n1929_ & ~new_n1940_;
  assign new_n1942_ = controlPi_67_5 & ~new_n1941_;
  assign new_n1943_ = ~new_n1907_ & ~new_n1942_;
  assign new_n1944_ = controlPi_67_0 & ~new_n1943_;
  assign new_n1945_ = ~controlPi_67_0 & new_n1943_;
  assign new_n1946_ = ~new_n1944_ & ~new_n1945_;
  assign new_n1947_ = ~new_n1861_ & ~new_n1946_;
  assign new_n1948_ = new_n1690_ & new_n1775_;
  assign new_n1949_ = new_n1947_ & ~new_n1948_;
  assign new_n1950_ = ~new_n1776_ & ~new_n1949_;
  assign new_n1951_ = ~controlPi_2_1 & ~n199_ntk1;
  assign new_n1952_ = controlPi_2_1 & ~n211_ntk1;
  assign new_n1953_ = ~new_n1951_ & ~new_n1952_;
  assign new_n1954_ = ~controlPi_2_2 & new_n1953_;
  assign new_n1955_ = ~controlPi_2_1 & ~n216_ntk1;
  assign new_n1956_ = controlPi_2_1 & ~n280_ntk1;
  assign new_n1957_ = ~new_n1955_ & ~new_n1956_;
  assign new_n1958_ = controlPi_2_2 & new_n1957_;
  assign new_n1959_ = ~new_n1954_ & ~new_n1958_;
  assign new_n1960_ = ~controlPi_2_3 & new_n1959_;
  assign new_n1961_ = ~controlPi_2_1 & ~n287_ntk1;
  assign new_n1962_ = controlPi_2_1 & ~n409_ntk1;
  assign new_n1963_ = ~new_n1961_ & ~new_n1962_;
  assign new_n1964_ = ~controlPi_2_2 & new_n1963_;
  assign new_n1965_ = ~controlPi_2_1 & ~n428_ntk1;
  assign new_n1966_ = controlPi_2_1 & ~n435_ntk1;
  assign new_n1967_ = ~new_n1965_ & ~new_n1966_;
  assign new_n1968_ = controlPi_2_2 & new_n1967_;
  assign new_n1969_ = ~new_n1964_ & ~new_n1968_;
  assign new_n1970_ = controlPi_2_3 & new_n1969_;
  assign new_n1971_ = ~new_n1960_ & ~new_n1970_;
  assign new_n1972_ = controlPi_2_4 & ~new_n1971_;
  assign new_n1973_ = ~controlPi_2_1 & ~n2_ntk1;
  assign new_n1974_ = controlPi_2_1 & ~n13_ntk1;
  assign new_n1975_ = ~new_n1973_ & ~new_n1974_;
  assign new_n1976_ = ~controlPi_2_2 & new_n1975_;
  assign new_n1977_ = ~controlPi_2_1 & ~n46_ntk1;
  assign new_n1978_ = controlPi_2_1 & ~n75_ntk1;
  assign new_n1979_ = ~new_n1977_ & ~new_n1978_;
  assign new_n1980_ = controlPi_2_2 & new_n1979_;
  assign new_n1981_ = ~new_n1976_ & ~new_n1980_;
  assign new_n1982_ = ~controlPi_2_3 & new_n1981_;
  assign new_n1983_ = ~controlPi_2_1 & ~n96_ntk1;
  assign new_n1984_ = controlPi_2_1 & ~n131_ntk1;
  assign new_n1985_ = ~new_n1983_ & ~new_n1984_;
  assign new_n1986_ = ~controlPi_2_2 & new_n1985_;
  assign new_n1987_ = ~controlPi_2_1 & ~n159_ntk1;
  assign new_n1988_ = controlPi_2_1 & ~n177_ntk1;
  assign new_n1989_ = ~new_n1987_ & ~new_n1988_;
  assign new_n1990_ = controlPi_2_2 & new_n1989_;
  assign new_n1991_ = ~new_n1986_ & ~new_n1990_;
  assign new_n1992_ = controlPi_2_3 & new_n1991_;
  assign new_n1993_ = ~new_n1982_ & ~new_n1992_;
  assign new_n1994_ = ~controlPi_2_4 & ~new_n1993_;
  assign new_n1995_ = ~new_n1972_ & ~new_n1994_;
  assign new_n1996_ = ~controlPi_2_5 & ~new_n1995_;
  assign new_n1997_ = controlPi_2_1 & n659_ntk1;
  assign new_n1998_ = ~controlPi_2_1 & n616_ntk1;
  assign new_n1999_ = ~new_n1997_ & ~new_n1998_;
  assign new_n2000_ = ~controlPi_2_2 & new_n1999_;
  assign new_n2001_ = controlPi_2_1 & n673_ntk1;
  assign new_n2002_ = ~controlPi_2_1 & n664_ntk1;
  assign new_n2003_ = ~new_n2001_ & ~new_n2002_;
  assign new_n2004_ = controlPi_2_2 & new_n2003_;
  assign new_n2005_ = ~new_n2000_ & ~new_n2004_;
  assign new_n2006_ = controlPi_2_4 & ~new_n2005_;
  assign new_n2007_ = controlPi_2_1 & n457_ntk1;
  assign new_n2008_ = ~controlPi_2_1 & n454_ntk1;
  assign new_n2009_ = ~new_n2007_ & ~new_n2008_;
  assign new_n2010_ = ~controlPi_2_2 & new_n2009_;
  assign new_n2011_ = controlPi_2_1 & n507_ntk1;
  assign new_n2012_ = ~controlPi_2_1 & n468_ntk1;
  assign new_n2013_ = ~new_n2011_ & ~new_n2012_;
  assign new_n2014_ = controlPi_2_2 & new_n2013_;
  assign new_n2015_ = ~new_n2010_ & ~new_n2014_;
  assign new_n2016_ = ~controlPi_2_4 & ~new_n2015_;
  assign new_n2017_ = ~new_n2006_ & ~new_n2016_;
  assign new_n2018_ = ~controlPi_2_3 & ~new_n2017_;
  assign new_n2019_ = controlPi_2_1 & n600_ntk1;
  assign new_n2020_ = ~controlPi_2_1 & n582_ntk1;
  assign new_n2021_ = ~new_n2019_ & ~new_n2020_;
  assign new_n2022_ = controlPi_2_2 & new_n2021_;
  assign new_n2023_ = controlPi_2_1 & n525_ntk1;
  assign new_n2024_ = ~controlPi_2_1 & n511_ntk1;
  assign new_n2025_ = ~new_n2023_ & ~new_n2024_;
  assign new_n2026_ = ~controlPi_2_2 & new_n2025_;
  assign new_n2027_ = ~new_n2022_ & ~new_n2026_;
  assign new_n2028_ = controlPi_2_3 & ~new_n2027_;
  assign new_n2029_ = ~controlPi_2_4 & new_n2028_;
  assign new_n2030_ = ~new_n2018_ & ~new_n2029_;
  assign new_n2031_ = controlPi_2_5 & ~new_n2030_;
  assign new_n2032_ = ~new_n1996_ & ~new_n2031_;
  assign new_n2033_ = controlPi_2_0 & ~new_n2032_;
  assign new_n2034_ = ~controlPi_2_0 & new_n2032_;
  assign new_n2035_ = ~new_n2033_ & ~new_n2034_;
  assign new_n2036_ = ~controlPi_74_1 & ~n199_ntk1;
  assign new_n2037_ = controlPi_74_1 & ~n211_ntk1;
  assign new_n2038_ = ~new_n2036_ & ~new_n2037_;
  assign new_n2039_ = ~controlPi_74_2 & new_n2038_;
  assign new_n2040_ = ~controlPi_74_1 & ~n216_ntk1;
  assign new_n2041_ = controlPi_74_1 & ~n280_ntk1;
  assign new_n2042_ = ~new_n2040_ & ~new_n2041_;
  assign new_n2043_ = controlPi_74_2 & new_n2042_;
  assign new_n2044_ = ~new_n2039_ & ~new_n2043_;
  assign new_n2045_ = ~controlPi_74_3 & new_n2044_;
  assign new_n2046_ = ~controlPi_74_1 & ~n287_ntk1;
  assign new_n2047_ = controlPi_74_1 & ~n409_ntk1;
  assign new_n2048_ = ~new_n2046_ & ~new_n2047_;
  assign new_n2049_ = ~controlPi_74_2 & new_n2048_;
  assign new_n2050_ = ~controlPi_74_1 & ~n428_ntk1;
  assign new_n2051_ = controlPi_74_1 & ~n435_ntk1;
  assign new_n2052_ = ~new_n2050_ & ~new_n2051_;
  assign new_n2053_ = controlPi_74_2 & new_n2052_;
  assign new_n2054_ = ~new_n2049_ & ~new_n2053_;
  assign new_n2055_ = controlPi_74_3 & new_n2054_;
  assign new_n2056_ = ~new_n2045_ & ~new_n2055_;
  assign new_n2057_ = controlPi_74_4 & ~new_n2056_;
  assign new_n2058_ = ~controlPi_74_1 & ~n2_ntk1;
  assign new_n2059_ = controlPi_74_1 & ~n13_ntk1;
  assign new_n2060_ = ~new_n2058_ & ~new_n2059_;
  assign new_n2061_ = ~controlPi_74_2 & new_n2060_;
  assign new_n2062_ = ~controlPi_74_1 & ~n46_ntk1;
  assign new_n2063_ = controlPi_74_1 & ~n75_ntk1;
  assign new_n2064_ = ~new_n2062_ & ~new_n2063_;
  assign new_n2065_ = controlPi_74_2 & new_n2064_;
  assign new_n2066_ = ~new_n2061_ & ~new_n2065_;
  assign new_n2067_ = ~controlPi_74_3 & new_n2066_;
  assign new_n2068_ = ~controlPi_74_1 & ~n96_ntk1;
  assign new_n2069_ = controlPi_74_1 & ~n131_ntk1;
  assign new_n2070_ = ~new_n2068_ & ~new_n2069_;
  assign new_n2071_ = ~controlPi_74_2 & new_n2070_;
  assign new_n2072_ = ~controlPi_74_1 & ~n159_ntk1;
  assign new_n2073_ = controlPi_74_1 & ~n177_ntk1;
  assign new_n2074_ = ~new_n2072_ & ~new_n2073_;
  assign new_n2075_ = controlPi_74_2 & new_n2074_;
  assign new_n2076_ = ~new_n2071_ & ~new_n2075_;
  assign new_n2077_ = controlPi_74_3 & new_n2076_;
  assign new_n2078_ = ~new_n2067_ & ~new_n2077_;
  assign new_n2079_ = ~controlPi_74_4 & ~new_n2078_;
  assign new_n2080_ = ~new_n2057_ & ~new_n2079_;
  assign new_n2081_ = ~controlPi_74_5 & ~new_n2080_;
  assign new_n2082_ = controlPi_74_1 & n659_ntk1;
  assign new_n2083_ = ~controlPi_74_1 & n616_ntk1;
  assign new_n2084_ = ~new_n2082_ & ~new_n2083_;
  assign new_n2085_ = ~controlPi_74_2 & new_n2084_;
  assign new_n2086_ = controlPi_74_1 & n673_ntk1;
  assign new_n2087_ = ~controlPi_74_1 & n664_ntk1;
  assign new_n2088_ = ~new_n2086_ & ~new_n2087_;
  assign new_n2089_ = controlPi_74_2 & new_n2088_;
  assign new_n2090_ = ~new_n2085_ & ~new_n2089_;
  assign new_n2091_ = controlPi_74_4 & ~new_n2090_;
  assign new_n2092_ = controlPi_74_1 & n457_ntk1;
  assign new_n2093_ = ~controlPi_74_1 & n454_ntk1;
  assign new_n2094_ = ~new_n2092_ & ~new_n2093_;
  assign new_n2095_ = ~controlPi_74_2 & new_n2094_;
  assign new_n2096_ = controlPi_74_1 & n507_ntk1;
  assign new_n2097_ = ~controlPi_74_1 & n468_ntk1;
  assign new_n2098_ = ~new_n2096_ & ~new_n2097_;
  assign new_n2099_ = controlPi_74_2 & new_n2098_;
  assign new_n2100_ = ~new_n2095_ & ~new_n2099_;
  assign new_n2101_ = ~controlPi_74_4 & ~new_n2100_;
  assign new_n2102_ = ~new_n2091_ & ~new_n2101_;
  assign new_n2103_ = ~controlPi_74_3 & ~new_n2102_;
  assign new_n2104_ = controlPi_74_1 & n600_ntk1;
  assign new_n2105_ = ~controlPi_74_1 & n582_ntk1;
  assign new_n2106_ = ~new_n2104_ & ~new_n2105_;
  assign new_n2107_ = controlPi_74_2 & new_n2106_;
  assign new_n2108_ = controlPi_74_1 & n525_ntk1;
  assign new_n2109_ = ~controlPi_74_1 & n511_ntk1;
  assign new_n2110_ = ~new_n2108_ & ~new_n2109_;
  assign new_n2111_ = ~controlPi_74_2 & new_n2110_;
  assign new_n2112_ = ~new_n2107_ & ~new_n2111_;
  assign new_n2113_ = controlPi_74_3 & ~new_n2112_;
  assign new_n2114_ = ~controlPi_74_4 & new_n2113_;
  assign new_n2115_ = ~new_n2103_ & ~new_n2114_;
  assign new_n2116_ = controlPi_74_5 & ~new_n2115_;
  assign new_n2117_ = ~new_n2081_ & ~new_n2116_;
  assign new_n2118_ = controlPi_74_0 & ~new_n2117_;
  assign new_n2119_ = ~controlPi_74_0 & new_n2117_;
  assign new_n2120_ = ~new_n2118_ & ~new_n2119_;
  assign new_n2121_ = new_n2035_ & new_n2120_;
  assign new_n2122_ = ~new_n2035_ & ~new_n2120_;
  assign new_n2123_ = ~new_n2121_ & ~new_n2122_;
  assign new_n2124_ = new_n1950_ & ~new_n2123_;
  assign new_n2125_ = ~new_n1950_ & new_n2123_;
  assign new_n2126_ = ~new_n2124_ & ~new_n2125_;
  assign new_n2127_ = ~new_n1605_ & ~new_n2126_;
  assign new_n2128_ = ~controlPi_36_1 & ~n349_ntk1;
  assign new_n2129_ = controlPi_36_1 & ~n368_ntk1;
  assign new_n2130_ = ~new_n2128_ & ~new_n2129_;
  assign new_n2131_ = controlPi_36_3 & ~new_n2130_;
  assign new_n2132_ = ~controlPi_36_1 & ~n85_ntk1;
  assign new_n2133_ = controlPi_36_1 & ~n93_ntk1;
  assign new_n2134_ = ~new_n2132_ & ~new_n2133_;
  assign new_n2135_ = ~controlPi_36_3 & ~new_n2134_;
  assign new_n2136_ = ~new_n2131_ & ~new_n2135_;
  assign new_n2137_ = ~controlPi_36_2 & ~new_n2136_;
  assign new_n2138_ = ~controlPi_36_1 & ~n206_ntk1;
  assign new_n2139_ = controlPi_36_1 & ~n266_ntk1;
  assign new_n2140_ = ~new_n2138_ & ~new_n2139_;
  assign new_n2141_ = controlPi_36_2 & ~new_n2140_;
  assign new_n2142_ = ~controlPi_36_3 & new_n2141_;
  assign new_n2143_ = ~new_n2137_ & ~new_n2142_;
  assign new_n2144_ = controlPi_36_0 & ~new_n2143_;
  assign new_n2145_ = ~controlPi_36_0 & new_n2143_;
  assign new_n2146_ = ~new_n2144_ & ~new_n2145_;
  assign new_n2147_ = ~controlPi_14_1 & ~n199_ntk1;
  assign new_n2148_ = controlPi_14_1 & ~n211_ntk1;
  assign new_n2149_ = ~new_n2147_ & ~new_n2148_;
  assign new_n2150_ = ~controlPi_14_2 & new_n2149_;
  assign new_n2151_ = ~controlPi_14_1 & ~n216_ntk1;
  assign new_n2152_ = controlPi_14_1 & ~n280_ntk1;
  assign new_n2153_ = ~new_n2151_ & ~new_n2152_;
  assign new_n2154_ = controlPi_14_2 & new_n2153_;
  assign new_n2155_ = ~new_n2150_ & ~new_n2154_;
  assign new_n2156_ = ~controlPi_14_3 & new_n2155_;
  assign new_n2157_ = ~controlPi_14_1 & ~n287_ntk1;
  assign new_n2158_ = controlPi_14_1 & ~n409_ntk1;
  assign new_n2159_ = ~new_n2157_ & ~new_n2158_;
  assign new_n2160_ = ~controlPi_14_2 & new_n2159_;
  assign new_n2161_ = ~controlPi_14_1 & ~n428_ntk1;
  assign new_n2162_ = controlPi_14_1 & ~n435_ntk1;
  assign new_n2163_ = ~new_n2161_ & ~new_n2162_;
  assign new_n2164_ = controlPi_14_2 & new_n2163_;
  assign new_n2165_ = ~new_n2160_ & ~new_n2164_;
  assign new_n2166_ = controlPi_14_3 & new_n2165_;
  assign new_n2167_ = ~new_n2156_ & ~new_n2166_;
  assign new_n2168_ = controlPi_14_4 & ~new_n2167_;
  assign new_n2169_ = ~controlPi_14_1 & ~n2_ntk1;
  assign new_n2170_ = controlPi_14_1 & ~n13_ntk1;
  assign new_n2171_ = ~new_n2169_ & ~new_n2170_;
  assign new_n2172_ = ~controlPi_14_2 & new_n2171_;
  assign new_n2173_ = ~controlPi_14_1 & ~n46_ntk1;
  assign new_n2174_ = controlPi_14_1 & ~n75_ntk1;
  assign new_n2175_ = ~new_n2173_ & ~new_n2174_;
  assign new_n2176_ = controlPi_14_2 & new_n2175_;
  assign new_n2177_ = ~new_n2172_ & ~new_n2176_;
  assign new_n2178_ = ~controlPi_14_3 & new_n2177_;
  assign new_n2179_ = ~controlPi_14_1 & ~n96_ntk1;
  assign new_n2180_ = controlPi_14_1 & ~n131_ntk1;
  assign new_n2181_ = ~new_n2179_ & ~new_n2180_;
  assign new_n2182_ = ~controlPi_14_2 & new_n2181_;
  assign new_n2183_ = ~controlPi_14_1 & ~n159_ntk1;
  assign new_n2184_ = controlPi_14_1 & ~n177_ntk1;
  assign new_n2185_ = ~new_n2183_ & ~new_n2184_;
  assign new_n2186_ = controlPi_14_2 & new_n2185_;
  assign new_n2187_ = ~new_n2182_ & ~new_n2186_;
  assign new_n2188_ = controlPi_14_3 & new_n2187_;
  assign new_n2189_ = ~new_n2178_ & ~new_n2188_;
  assign new_n2190_ = ~controlPi_14_4 & ~new_n2189_;
  assign new_n2191_ = ~new_n2168_ & ~new_n2190_;
  assign new_n2192_ = ~controlPi_14_5 & ~new_n2191_;
  assign new_n2193_ = controlPi_14_1 & n659_ntk1;
  assign new_n2194_ = ~controlPi_14_1 & n616_ntk1;
  assign new_n2195_ = ~new_n2193_ & ~new_n2194_;
  assign new_n2196_ = ~controlPi_14_2 & new_n2195_;
  assign new_n2197_ = controlPi_14_1 & n673_ntk1;
  assign new_n2198_ = ~controlPi_14_1 & n664_ntk1;
  assign new_n2199_ = ~new_n2197_ & ~new_n2198_;
  assign new_n2200_ = controlPi_14_2 & new_n2199_;
  assign new_n2201_ = ~new_n2196_ & ~new_n2200_;
  assign new_n2202_ = controlPi_14_4 & ~new_n2201_;
  assign new_n2203_ = controlPi_14_1 & n457_ntk1;
  assign new_n2204_ = ~controlPi_14_1 & n454_ntk1;
  assign new_n2205_ = ~new_n2203_ & ~new_n2204_;
  assign new_n2206_ = ~controlPi_14_2 & new_n2205_;
  assign new_n2207_ = controlPi_14_1 & n507_ntk1;
  assign new_n2208_ = ~controlPi_14_1 & n468_ntk1;
  assign new_n2209_ = ~new_n2207_ & ~new_n2208_;
  assign new_n2210_ = controlPi_14_2 & new_n2209_;
  assign new_n2211_ = ~new_n2206_ & ~new_n2210_;
  assign new_n2212_ = ~controlPi_14_4 & ~new_n2211_;
  assign new_n2213_ = ~new_n2202_ & ~new_n2212_;
  assign new_n2214_ = ~controlPi_14_3 & ~new_n2213_;
  assign new_n2215_ = controlPi_14_1 & n600_ntk1;
  assign new_n2216_ = ~controlPi_14_1 & n582_ntk1;
  assign new_n2217_ = ~new_n2215_ & ~new_n2216_;
  assign new_n2218_ = controlPi_14_2 & new_n2217_;
  assign new_n2219_ = controlPi_14_1 & n525_ntk1;
  assign new_n2220_ = ~controlPi_14_1 & n511_ntk1;
  assign new_n2221_ = ~new_n2219_ & ~new_n2220_;
  assign new_n2222_ = ~controlPi_14_2 & new_n2221_;
  assign new_n2223_ = ~new_n2218_ & ~new_n2222_;
  assign new_n2224_ = controlPi_14_3 & ~new_n2223_;
  assign new_n2225_ = ~controlPi_14_4 & new_n2224_;
  assign new_n2226_ = ~new_n2214_ & ~new_n2225_;
  assign new_n2227_ = controlPi_14_5 & ~new_n2226_;
  assign new_n2228_ = ~new_n2192_ & ~new_n2227_;
  assign new_n2229_ = controlPi_14_0 & ~new_n2228_;
  assign new_n2230_ = ~controlPi_14_0 & new_n2228_;
  assign new_n2231_ = ~new_n2229_ & ~new_n2230_;
  assign new_n2232_ = ~new_n1775_ & ~new_n2231_;
  assign new_n2233_ = ~controlPi_66_1 & ~n199_ntk1;
  assign new_n2234_ = controlPi_66_1 & ~n211_ntk1;
  assign new_n2235_ = ~new_n2233_ & ~new_n2234_;
  assign new_n2236_ = ~controlPi_66_2 & new_n2235_;
  assign new_n2237_ = ~controlPi_66_1 & ~n216_ntk1;
  assign new_n2238_ = controlPi_66_1 & ~n280_ntk1;
  assign new_n2239_ = ~new_n2237_ & ~new_n2238_;
  assign new_n2240_ = controlPi_66_2 & new_n2239_;
  assign new_n2241_ = ~new_n2236_ & ~new_n2240_;
  assign new_n2242_ = ~controlPi_66_3 & new_n2241_;
  assign new_n2243_ = ~controlPi_66_1 & ~n287_ntk1;
  assign new_n2244_ = controlPi_66_1 & ~n409_ntk1;
  assign new_n2245_ = ~new_n2243_ & ~new_n2244_;
  assign new_n2246_ = ~controlPi_66_2 & new_n2245_;
  assign new_n2247_ = ~controlPi_66_1 & ~n428_ntk1;
  assign new_n2248_ = controlPi_66_1 & ~n435_ntk1;
  assign new_n2249_ = ~new_n2247_ & ~new_n2248_;
  assign new_n2250_ = controlPi_66_2 & new_n2249_;
  assign new_n2251_ = ~new_n2246_ & ~new_n2250_;
  assign new_n2252_ = controlPi_66_3 & new_n2251_;
  assign new_n2253_ = ~new_n2242_ & ~new_n2252_;
  assign new_n2254_ = controlPi_66_4 & ~new_n2253_;
  assign new_n2255_ = ~controlPi_66_1 & ~n2_ntk1;
  assign new_n2256_ = controlPi_66_1 & ~n13_ntk1;
  assign new_n2257_ = ~new_n2255_ & ~new_n2256_;
  assign new_n2258_ = ~controlPi_66_2 & new_n2257_;
  assign new_n2259_ = ~controlPi_66_1 & ~n46_ntk1;
  assign new_n2260_ = controlPi_66_1 & ~n75_ntk1;
  assign new_n2261_ = ~new_n2259_ & ~new_n2260_;
  assign new_n2262_ = controlPi_66_2 & new_n2261_;
  assign new_n2263_ = ~new_n2258_ & ~new_n2262_;
  assign new_n2264_ = ~controlPi_66_3 & new_n2263_;
  assign new_n2265_ = ~controlPi_66_1 & ~n96_ntk1;
  assign new_n2266_ = controlPi_66_1 & ~n131_ntk1;
  assign new_n2267_ = ~new_n2265_ & ~new_n2266_;
  assign new_n2268_ = ~controlPi_66_2 & new_n2267_;
  assign new_n2269_ = ~controlPi_66_1 & ~n159_ntk1;
  assign new_n2270_ = controlPi_66_1 & ~n177_ntk1;
  assign new_n2271_ = ~new_n2269_ & ~new_n2270_;
  assign new_n2272_ = controlPi_66_2 & new_n2271_;
  assign new_n2273_ = ~new_n2268_ & ~new_n2272_;
  assign new_n2274_ = controlPi_66_3 & new_n2273_;
  assign new_n2275_ = ~new_n2264_ & ~new_n2274_;
  assign new_n2276_ = ~controlPi_66_4 & ~new_n2275_;
  assign new_n2277_ = ~new_n2254_ & ~new_n2276_;
  assign new_n2278_ = ~controlPi_66_5 & ~new_n2277_;
  assign new_n2279_ = controlPi_66_1 & n659_ntk1;
  assign new_n2280_ = ~controlPi_66_1 & n616_ntk1;
  assign new_n2281_ = ~new_n2279_ & ~new_n2280_;
  assign new_n2282_ = ~controlPi_66_2 & new_n2281_;
  assign new_n2283_ = controlPi_66_1 & n673_ntk1;
  assign new_n2284_ = ~controlPi_66_1 & n664_ntk1;
  assign new_n2285_ = ~new_n2283_ & ~new_n2284_;
  assign new_n2286_ = controlPi_66_2 & new_n2285_;
  assign new_n2287_ = ~new_n2282_ & ~new_n2286_;
  assign new_n2288_ = controlPi_66_4 & ~new_n2287_;
  assign new_n2289_ = controlPi_66_1 & n457_ntk1;
  assign new_n2290_ = ~controlPi_66_1 & n454_ntk1;
  assign new_n2291_ = ~new_n2289_ & ~new_n2290_;
  assign new_n2292_ = ~controlPi_66_2 & new_n2291_;
  assign new_n2293_ = controlPi_66_1 & n507_ntk1;
  assign new_n2294_ = ~controlPi_66_1 & n468_ntk1;
  assign new_n2295_ = ~new_n2293_ & ~new_n2294_;
  assign new_n2296_ = controlPi_66_2 & new_n2295_;
  assign new_n2297_ = ~new_n2292_ & ~new_n2296_;
  assign new_n2298_ = ~controlPi_66_4 & ~new_n2297_;
  assign new_n2299_ = ~new_n2288_ & ~new_n2298_;
  assign new_n2300_ = ~controlPi_66_3 & ~new_n2299_;
  assign new_n2301_ = controlPi_66_1 & n600_ntk1;
  assign new_n2302_ = ~controlPi_66_1 & n582_ntk1;
  assign new_n2303_ = ~new_n2301_ & ~new_n2302_;
  assign new_n2304_ = controlPi_66_2 & new_n2303_;
  assign new_n2305_ = controlPi_66_1 & n525_ntk1;
  assign new_n2306_ = ~controlPi_66_1 & n511_ntk1;
  assign new_n2307_ = ~new_n2305_ & ~new_n2306_;
  assign new_n2308_ = ~controlPi_66_2 & new_n2307_;
  assign new_n2309_ = ~new_n2304_ & ~new_n2308_;
  assign new_n2310_ = controlPi_66_3 & ~new_n2309_;
  assign new_n2311_ = ~controlPi_66_4 & new_n2310_;
  assign new_n2312_ = ~new_n2300_ & ~new_n2311_;
  assign new_n2313_ = controlPi_66_5 & ~new_n2312_;
  assign new_n2314_ = ~new_n2278_ & ~new_n2313_;
  assign new_n2315_ = controlPi_66_0 & ~new_n2314_;
  assign new_n2316_ = ~controlPi_66_0 & new_n2314_;
  assign new_n2317_ = ~new_n2315_ & ~new_n2316_;
  assign new_n2318_ = ~new_n1946_ & ~new_n2317_;
  assign new_n2319_ = new_n1775_ & new_n2231_;
  assign new_n2320_ = new_n2318_ & ~new_n2319_;
  assign new_n2321_ = ~new_n2232_ & ~new_n2320_;
  assign new_n2322_ = ~controlPi_84_1 & ~n199_ntk1;
  assign new_n2323_ = controlPi_84_1 & ~n211_ntk1;
  assign new_n2324_ = ~new_n2322_ & ~new_n2323_;
  assign new_n2325_ = ~controlPi_84_2 & new_n2324_;
  assign new_n2326_ = ~controlPi_84_1 & ~n216_ntk1;
  assign new_n2327_ = controlPi_84_1 & ~n280_ntk1;
  assign new_n2328_ = ~new_n2326_ & ~new_n2327_;
  assign new_n2329_ = controlPi_84_2 & new_n2328_;
  assign new_n2330_ = ~new_n2325_ & ~new_n2329_;
  assign new_n2331_ = ~controlPi_84_3 & new_n2330_;
  assign new_n2332_ = ~controlPi_84_1 & ~n287_ntk1;
  assign new_n2333_ = controlPi_84_1 & ~n409_ntk1;
  assign new_n2334_ = ~new_n2332_ & ~new_n2333_;
  assign new_n2335_ = ~controlPi_84_2 & new_n2334_;
  assign new_n2336_ = ~controlPi_84_1 & ~n428_ntk1;
  assign new_n2337_ = controlPi_84_1 & ~n435_ntk1;
  assign new_n2338_ = ~new_n2336_ & ~new_n2337_;
  assign new_n2339_ = controlPi_84_2 & new_n2338_;
  assign new_n2340_ = ~new_n2335_ & ~new_n2339_;
  assign new_n2341_ = controlPi_84_3 & new_n2340_;
  assign new_n2342_ = ~new_n2331_ & ~new_n2341_;
  assign new_n2343_ = controlPi_84_4 & ~new_n2342_;
  assign new_n2344_ = ~controlPi_84_1 & ~n2_ntk1;
  assign new_n2345_ = controlPi_84_1 & ~n13_ntk1;
  assign new_n2346_ = ~new_n2344_ & ~new_n2345_;
  assign new_n2347_ = ~controlPi_84_2 & new_n2346_;
  assign new_n2348_ = ~controlPi_84_1 & ~n46_ntk1;
  assign new_n2349_ = controlPi_84_1 & ~n75_ntk1;
  assign new_n2350_ = ~new_n2348_ & ~new_n2349_;
  assign new_n2351_ = controlPi_84_2 & new_n2350_;
  assign new_n2352_ = ~new_n2347_ & ~new_n2351_;
  assign new_n2353_ = ~controlPi_84_3 & new_n2352_;
  assign new_n2354_ = ~controlPi_84_1 & ~n96_ntk1;
  assign new_n2355_ = controlPi_84_1 & ~n131_ntk1;
  assign new_n2356_ = ~new_n2354_ & ~new_n2355_;
  assign new_n2357_ = ~controlPi_84_2 & new_n2356_;
  assign new_n2358_ = ~controlPi_84_1 & ~n159_ntk1;
  assign new_n2359_ = controlPi_84_1 & ~n177_ntk1;
  assign new_n2360_ = ~new_n2358_ & ~new_n2359_;
  assign new_n2361_ = controlPi_84_2 & new_n2360_;
  assign new_n2362_ = ~new_n2357_ & ~new_n2361_;
  assign new_n2363_ = controlPi_84_3 & new_n2362_;
  assign new_n2364_ = ~new_n2353_ & ~new_n2363_;
  assign new_n2365_ = ~controlPi_84_4 & ~new_n2364_;
  assign new_n2366_ = ~new_n2343_ & ~new_n2365_;
  assign new_n2367_ = ~controlPi_84_5 & ~new_n2366_;
  assign new_n2368_ = controlPi_84_1 & n659_ntk1;
  assign new_n2369_ = ~controlPi_84_1 & n616_ntk1;
  assign new_n2370_ = ~new_n2368_ & ~new_n2369_;
  assign new_n2371_ = ~controlPi_84_2 & new_n2370_;
  assign new_n2372_ = controlPi_84_1 & n673_ntk1;
  assign new_n2373_ = ~controlPi_84_1 & n664_ntk1;
  assign new_n2374_ = ~new_n2372_ & ~new_n2373_;
  assign new_n2375_ = controlPi_84_2 & new_n2374_;
  assign new_n2376_ = ~new_n2371_ & ~new_n2375_;
  assign new_n2377_ = controlPi_84_4 & ~new_n2376_;
  assign new_n2378_ = controlPi_84_1 & n457_ntk1;
  assign new_n2379_ = ~controlPi_84_1 & n454_ntk1;
  assign new_n2380_ = ~new_n2378_ & ~new_n2379_;
  assign new_n2381_ = ~controlPi_84_2 & new_n2380_;
  assign new_n2382_ = controlPi_84_1 & n507_ntk1;
  assign new_n2383_ = ~controlPi_84_1 & n468_ntk1;
  assign new_n2384_ = ~new_n2382_ & ~new_n2383_;
  assign new_n2385_ = controlPi_84_2 & new_n2384_;
  assign new_n2386_ = ~new_n2381_ & ~new_n2385_;
  assign new_n2387_ = ~controlPi_84_4 & ~new_n2386_;
  assign new_n2388_ = ~new_n2377_ & ~new_n2387_;
  assign new_n2389_ = ~controlPi_84_3 & ~new_n2388_;
  assign new_n2390_ = controlPi_84_1 & n600_ntk1;
  assign new_n2391_ = ~controlPi_84_1 & n582_ntk1;
  assign new_n2392_ = ~new_n2390_ & ~new_n2391_;
  assign new_n2393_ = controlPi_84_2 & new_n2392_;
  assign new_n2394_ = controlPi_84_1 & n525_ntk1;
  assign new_n2395_ = ~controlPi_84_1 & n511_ntk1;
  assign new_n2396_ = ~new_n2394_ & ~new_n2395_;
  assign new_n2397_ = ~controlPi_84_2 & new_n2396_;
  assign new_n2398_ = ~new_n2393_ & ~new_n2397_;
  assign new_n2399_ = controlPi_84_3 & ~new_n2398_;
  assign new_n2400_ = ~controlPi_84_4 & new_n2399_;
  assign new_n2401_ = ~new_n2389_ & ~new_n2400_;
  assign new_n2402_ = controlPi_84_5 & ~new_n2401_;
  assign new_n2403_ = ~new_n2367_ & ~new_n2402_;
  assign new_n2404_ = controlPi_84_0 & ~new_n2403_;
  assign new_n2405_ = ~controlPi_84_0 & new_n2403_;
  assign new_n2406_ = ~new_n2404_ & ~new_n2405_;
  assign new_n2407_ = new_n2035_ & new_n2406_;
  assign new_n2408_ = ~new_n2035_ & ~new_n2406_;
  assign new_n2409_ = ~new_n2407_ & ~new_n2408_;
  assign new_n2410_ = new_n2321_ & ~new_n2409_;
  assign new_n2411_ = ~new_n2321_ & new_n2409_;
  assign new_n2412_ = ~new_n2410_ & ~new_n2411_;
  assign new_n2413_ = ~new_n2146_ & ~new_n2412_;
  assign new_n2414_ = ~controlPi_12_1 & ~n349_ntk1;
  assign new_n2415_ = controlPi_12_1 & ~n368_ntk1;
  assign new_n2416_ = ~new_n2414_ & ~new_n2415_;
  assign new_n2417_ = controlPi_12_3 & ~new_n2416_;
  assign new_n2418_ = ~controlPi_12_1 & ~n85_ntk1;
  assign new_n2419_ = controlPi_12_1 & ~n93_ntk1;
  assign new_n2420_ = ~new_n2418_ & ~new_n2419_;
  assign new_n2421_ = ~controlPi_12_3 & ~new_n2420_;
  assign new_n2422_ = ~new_n2417_ & ~new_n2421_;
  assign new_n2423_ = ~controlPi_12_2 & ~new_n2422_;
  assign new_n2424_ = ~controlPi_12_1 & ~n206_ntk1;
  assign new_n2425_ = controlPi_12_1 & ~n266_ntk1;
  assign new_n2426_ = ~new_n2424_ & ~new_n2425_;
  assign new_n2427_ = controlPi_12_2 & ~new_n2426_;
  assign new_n2428_ = ~controlPi_12_3 & new_n2427_;
  assign new_n2429_ = ~new_n2423_ & ~new_n2428_;
  assign new_n2430_ = controlPi_12_0 & ~new_n2429_;
  assign new_n2431_ = ~controlPi_12_0 & new_n2429_;
  assign new_n2432_ = ~new_n2430_ & ~new_n2431_;
  assign new_n2433_ = ~controlPi_52_1 & ~n199_ntk1;
  assign new_n2434_ = controlPi_52_1 & ~n211_ntk1;
  assign new_n2435_ = ~new_n2433_ & ~new_n2434_;
  assign new_n2436_ = ~controlPi_52_2 & new_n2435_;
  assign new_n2437_ = ~controlPi_52_1 & ~n216_ntk1;
  assign new_n2438_ = controlPi_52_1 & ~n280_ntk1;
  assign new_n2439_ = ~new_n2437_ & ~new_n2438_;
  assign new_n2440_ = controlPi_52_2 & new_n2439_;
  assign new_n2441_ = ~new_n2436_ & ~new_n2440_;
  assign new_n2442_ = ~controlPi_52_3 & new_n2441_;
  assign new_n2443_ = ~controlPi_52_1 & ~n287_ntk1;
  assign new_n2444_ = controlPi_52_1 & ~n409_ntk1;
  assign new_n2445_ = ~new_n2443_ & ~new_n2444_;
  assign new_n2446_ = ~controlPi_52_2 & new_n2445_;
  assign new_n2447_ = ~controlPi_52_1 & ~n428_ntk1;
  assign new_n2448_ = controlPi_52_1 & ~n435_ntk1;
  assign new_n2449_ = ~new_n2447_ & ~new_n2448_;
  assign new_n2450_ = controlPi_52_2 & new_n2449_;
  assign new_n2451_ = ~new_n2446_ & ~new_n2450_;
  assign new_n2452_ = controlPi_52_3 & new_n2451_;
  assign new_n2453_ = ~new_n2442_ & ~new_n2452_;
  assign new_n2454_ = controlPi_52_4 & ~new_n2453_;
  assign new_n2455_ = ~controlPi_52_1 & ~n2_ntk1;
  assign new_n2456_ = controlPi_52_1 & ~n13_ntk1;
  assign new_n2457_ = ~new_n2455_ & ~new_n2456_;
  assign new_n2458_ = ~controlPi_52_2 & new_n2457_;
  assign new_n2459_ = ~controlPi_52_1 & ~n46_ntk1;
  assign new_n2460_ = controlPi_52_1 & ~n75_ntk1;
  assign new_n2461_ = ~new_n2459_ & ~new_n2460_;
  assign new_n2462_ = controlPi_52_2 & new_n2461_;
  assign new_n2463_ = ~new_n2458_ & ~new_n2462_;
  assign new_n2464_ = ~controlPi_52_3 & new_n2463_;
  assign new_n2465_ = ~controlPi_52_1 & ~n96_ntk1;
  assign new_n2466_ = controlPi_52_1 & ~n131_ntk1;
  assign new_n2467_ = ~new_n2465_ & ~new_n2466_;
  assign new_n2468_ = ~controlPi_52_2 & new_n2467_;
  assign new_n2469_ = ~controlPi_52_1 & ~n159_ntk1;
  assign new_n2470_ = controlPi_52_1 & ~n177_ntk1;
  assign new_n2471_ = ~new_n2469_ & ~new_n2470_;
  assign new_n2472_ = controlPi_52_2 & new_n2471_;
  assign new_n2473_ = ~new_n2468_ & ~new_n2472_;
  assign new_n2474_ = controlPi_52_3 & new_n2473_;
  assign new_n2475_ = ~new_n2464_ & ~new_n2474_;
  assign new_n2476_ = ~controlPi_52_4 & ~new_n2475_;
  assign new_n2477_ = ~new_n2454_ & ~new_n2476_;
  assign new_n2478_ = ~controlPi_52_5 & ~new_n2477_;
  assign new_n2479_ = controlPi_52_1 & n659_ntk1;
  assign new_n2480_ = ~controlPi_52_1 & n616_ntk1;
  assign new_n2481_ = ~new_n2479_ & ~new_n2480_;
  assign new_n2482_ = ~controlPi_52_2 & new_n2481_;
  assign new_n2483_ = controlPi_52_1 & n673_ntk1;
  assign new_n2484_ = ~controlPi_52_1 & n664_ntk1;
  assign new_n2485_ = ~new_n2483_ & ~new_n2484_;
  assign new_n2486_ = controlPi_52_2 & new_n2485_;
  assign new_n2487_ = ~new_n2482_ & ~new_n2486_;
  assign new_n2488_ = controlPi_52_4 & ~new_n2487_;
  assign new_n2489_ = controlPi_52_1 & n457_ntk1;
  assign new_n2490_ = ~controlPi_52_1 & n454_ntk1;
  assign new_n2491_ = ~new_n2489_ & ~new_n2490_;
  assign new_n2492_ = ~controlPi_52_2 & new_n2491_;
  assign new_n2493_ = controlPi_52_1 & n507_ntk1;
  assign new_n2494_ = ~controlPi_52_1 & n468_ntk1;
  assign new_n2495_ = ~new_n2493_ & ~new_n2494_;
  assign new_n2496_ = controlPi_52_2 & new_n2495_;
  assign new_n2497_ = ~new_n2492_ & ~new_n2496_;
  assign new_n2498_ = ~controlPi_52_4 & ~new_n2497_;
  assign new_n2499_ = ~new_n2488_ & ~new_n2498_;
  assign new_n2500_ = ~controlPi_52_3 & ~new_n2499_;
  assign new_n2501_ = controlPi_52_1 & n600_ntk1;
  assign new_n2502_ = ~controlPi_52_1 & n582_ntk1;
  assign new_n2503_ = ~new_n2501_ & ~new_n2502_;
  assign new_n2504_ = controlPi_52_2 & new_n2503_;
  assign new_n2505_ = controlPi_52_1 & n525_ntk1;
  assign new_n2506_ = ~controlPi_52_1 & n511_ntk1;
  assign new_n2507_ = ~new_n2505_ & ~new_n2506_;
  assign new_n2508_ = ~controlPi_52_2 & new_n2507_;
  assign new_n2509_ = ~new_n2504_ & ~new_n2508_;
  assign new_n2510_ = controlPi_52_3 & ~new_n2509_;
  assign new_n2511_ = ~controlPi_52_4 & new_n2510_;
  assign new_n2512_ = ~new_n2500_ & ~new_n2511_;
  assign new_n2513_ = controlPi_52_5 & ~new_n2512_;
  assign new_n2514_ = ~new_n2478_ & ~new_n2513_;
  assign new_n2515_ = controlPi_52_0 & ~new_n2514_;
  assign new_n2516_ = ~controlPi_52_0 & new_n2514_;
  assign new_n2517_ = ~new_n2515_ & ~new_n2516_;
  assign new_n2518_ = new_n2432_ & new_n2517_;
  assign new_n2519_ = ~controlPi_80_1 & ~n199_ntk1;
  assign new_n2520_ = controlPi_80_1 & ~n211_ntk1;
  assign new_n2521_ = ~new_n2519_ & ~new_n2520_;
  assign new_n2522_ = ~controlPi_80_2 & new_n2521_;
  assign new_n2523_ = ~controlPi_80_1 & ~n216_ntk1;
  assign new_n2524_ = controlPi_80_1 & ~n280_ntk1;
  assign new_n2525_ = ~new_n2523_ & ~new_n2524_;
  assign new_n2526_ = controlPi_80_2 & new_n2525_;
  assign new_n2527_ = ~new_n2522_ & ~new_n2526_;
  assign new_n2528_ = ~controlPi_80_3 & new_n2527_;
  assign new_n2529_ = ~controlPi_80_1 & ~n287_ntk1;
  assign new_n2530_ = controlPi_80_1 & ~n409_ntk1;
  assign new_n2531_ = ~new_n2529_ & ~new_n2530_;
  assign new_n2532_ = ~controlPi_80_2 & new_n2531_;
  assign new_n2533_ = ~controlPi_80_1 & ~n428_ntk1;
  assign new_n2534_ = controlPi_80_1 & ~n435_ntk1;
  assign new_n2535_ = ~new_n2533_ & ~new_n2534_;
  assign new_n2536_ = controlPi_80_2 & new_n2535_;
  assign new_n2537_ = ~new_n2532_ & ~new_n2536_;
  assign new_n2538_ = controlPi_80_3 & new_n2537_;
  assign new_n2539_ = ~new_n2528_ & ~new_n2538_;
  assign new_n2540_ = controlPi_80_4 & ~new_n2539_;
  assign new_n2541_ = ~controlPi_80_1 & ~n2_ntk1;
  assign new_n2542_ = controlPi_80_1 & ~n13_ntk1;
  assign new_n2543_ = ~new_n2541_ & ~new_n2542_;
  assign new_n2544_ = ~controlPi_80_2 & new_n2543_;
  assign new_n2545_ = ~controlPi_80_1 & ~n46_ntk1;
  assign new_n2546_ = controlPi_80_1 & ~n75_ntk1;
  assign new_n2547_ = ~new_n2545_ & ~new_n2546_;
  assign new_n2548_ = controlPi_80_2 & new_n2547_;
  assign new_n2549_ = ~new_n2544_ & ~new_n2548_;
  assign new_n2550_ = ~controlPi_80_3 & new_n2549_;
  assign new_n2551_ = ~controlPi_80_1 & ~n96_ntk1;
  assign new_n2552_ = controlPi_80_1 & ~n131_ntk1;
  assign new_n2553_ = ~new_n2551_ & ~new_n2552_;
  assign new_n2554_ = ~controlPi_80_2 & new_n2553_;
  assign new_n2555_ = ~controlPi_80_1 & ~n159_ntk1;
  assign new_n2556_ = controlPi_80_1 & ~n177_ntk1;
  assign new_n2557_ = ~new_n2555_ & ~new_n2556_;
  assign new_n2558_ = controlPi_80_2 & new_n2557_;
  assign new_n2559_ = ~new_n2554_ & ~new_n2558_;
  assign new_n2560_ = controlPi_80_3 & new_n2559_;
  assign new_n2561_ = ~new_n2550_ & ~new_n2560_;
  assign new_n2562_ = ~controlPi_80_4 & ~new_n2561_;
  assign new_n2563_ = ~new_n2540_ & ~new_n2562_;
  assign new_n2564_ = ~controlPi_80_5 & ~new_n2563_;
  assign new_n2565_ = controlPi_80_1 & n659_ntk1;
  assign new_n2566_ = ~controlPi_80_1 & n616_ntk1;
  assign new_n2567_ = ~new_n2565_ & ~new_n2566_;
  assign new_n2568_ = ~controlPi_80_2 & new_n2567_;
  assign new_n2569_ = controlPi_80_1 & n673_ntk1;
  assign new_n2570_ = ~controlPi_80_1 & n664_ntk1;
  assign new_n2571_ = ~new_n2569_ & ~new_n2570_;
  assign new_n2572_ = controlPi_80_2 & new_n2571_;
  assign new_n2573_ = ~new_n2568_ & ~new_n2572_;
  assign new_n2574_ = controlPi_80_4 & ~new_n2573_;
  assign new_n2575_ = controlPi_80_1 & n457_ntk1;
  assign new_n2576_ = ~controlPi_80_1 & n454_ntk1;
  assign new_n2577_ = ~new_n2575_ & ~new_n2576_;
  assign new_n2578_ = ~controlPi_80_2 & new_n2577_;
  assign new_n2579_ = controlPi_80_1 & n507_ntk1;
  assign new_n2580_ = ~controlPi_80_1 & n468_ntk1;
  assign new_n2581_ = ~new_n2579_ & ~new_n2580_;
  assign new_n2582_ = controlPi_80_2 & new_n2581_;
  assign new_n2583_ = ~new_n2578_ & ~new_n2582_;
  assign new_n2584_ = ~controlPi_80_4 & ~new_n2583_;
  assign new_n2585_ = ~new_n2574_ & ~new_n2584_;
  assign new_n2586_ = ~controlPi_80_3 & ~new_n2585_;
  assign new_n2587_ = controlPi_80_1 & n600_ntk1;
  assign new_n2588_ = ~controlPi_80_1 & n582_ntk1;
  assign new_n2589_ = ~new_n2587_ & ~new_n2588_;
  assign new_n2590_ = controlPi_80_2 & new_n2589_;
  assign new_n2591_ = controlPi_80_1 & n525_ntk1;
  assign new_n2592_ = ~controlPi_80_1 & n511_ntk1;
  assign new_n2593_ = ~new_n2591_ & ~new_n2592_;
  assign new_n2594_ = ~controlPi_80_2 & new_n2593_;
  assign new_n2595_ = ~new_n2590_ & ~new_n2594_;
  assign new_n2596_ = controlPi_80_3 & ~new_n2595_;
  assign new_n2597_ = ~controlPi_80_4 & new_n2596_;
  assign new_n2598_ = ~new_n2586_ & ~new_n2597_;
  assign new_n2599_ = controlPi_80_5 & ~new_n2598_;
  assign new_n2600_ = ~new_n2564_ & ~new_n2599_;
  assign new_n2601_ = controlPi_80_0 & ~new_n2600_;
  assign new_n2602_ = ~controlPi_80_0 & new_n2600_;
  assign new_n2603_ = ~new_n2601_ & ~new_n2602_;
  assign new_n2604_ = ~new_n1775_ & ~new_n2603_;
  assign new_n2605_ = ~controlPi_13_1 & ~n199_ntk1;
  assign new_n2606_ = controlPi_13_1 & ~n211_ntk1;
  assign new_n2607_ = ~new_n2605_ & ~new_n2606_;
  assign new_n2608_ = ~controlPi_13_2 & new_n2607_;
  assign new_n2609_ = ~controlPi_13_1 & ~n216_ntk1;
  assign new_n2610_ = controlPi_13_1 & ~n280_ntk1;
  assign new_n2611_ = ~new_n2609_ & ~new_n2610_;
  assign new_n2612_ = controlPi_13_2 & new_n2611_;
  assign new_n2613_ = ~new_n2608_ & ~new_n2612_;
  assign new_n2614_ = ~controlPi_13_3 & new_n2613_;
  assign new_n2615_ = ~controlPi_13_1 & ~n287_ntk1;
  assign new_n2616_ = controlPi_13_1 & ~n409_ntk1;
  assign new_n2617_ = ~new_n2615_ & ~new_n2616_;
  assign new_n2618_ = ~controlPi_13_2 & new_n2617_;
  assign new_n2619_ = ~controlPi_13_1 & ~n428_ntk1;
  assign new_n2620_ = controlPi_13_1 & ~n435_ntk1;
  assign new_n2621_ = ~new_n2619_ & ~new_n2620_;
  assign new_n2622_ = controlPi_13_2 & new_n2621_;
  assign new_n2623_ = ~new_n2618_ & ~new_n2622_;
  assign new_n2624_ = controlPi_13_3 & new_n2623_;
  assign new_n2625_ = ~new_n2614_ & ~new_n2624_;
  assign new_n2626_ = controlPi_13_4 & ~new_n2625_;
  assign new_n2627_ = ~controlPi_13_1 & ~n2_ntk1;
  assign new_n2628_ = controlPi_13_1 & ~n13_ntk1;
  assign new_n2629_ = ~new_n2627_ & ~new_n2628_;
  assign new_n2630_ = ~controlPi_13_2 & new_n2629_;
  assign new_n2631_ = ~controlPi_13_1 & ~n46_ntk1;
  assign new_n2632_ = controlPi_13_1 & ~n75_ntk1;
  assign new_n2633_ = ~new_n2631_ & ~new_n2632_;
  assign new_n2634_ = controlPi_13_2 & new_n2633_;
  assign new_n2635_ = ~new_n2630_ & ~new_n2634_;
  assign new_n2636_ = ~controlPi_13_3 & new_n2635_;
  assign new_n2637_ = ~controlPi_13_1 & ~n96_ntk1;
  assign new_n2638_ = controlPi_13_1 & ~n131_ntk1;
  assign new_n2639_ = ~new_n2637_ & ~new_n2638_;
  assign new_n2640_ = ~controlPi_13_2 & new_n2639_;
  assign new_n2641_ = ~controlPi_13_1 & ~n159_ntk1;
  assign new_n2642_ = controlPi_13_1 & ~n177_ntk1;
  assign new_n2643_ = ~new_n2641_ & ~new_n2642_;
  assign new_n2644_ = controlPi_13_2 & new_n2643_;
  assign new_n2645_ = ~new_n2640_ & ~new_n2644_;
  assign new_n2646_ = controlPi_13_3 & new_n2645_;
  assign new_n2647_ = ~new_n2636_ & ~new_n2646_;
  assign new_n2648_ = ~controlPi_13_4 & ~new_n2647_;
  assign new_n2649_ = ~new_n2626_ & ~new_n2648_;
  assign new_n2650_ = ~controlPi_13_5 & ~new_n2649_;
  assign new_n2651_ = controlPi_13_1 & n659_ntk1;
  assign new_n2652_ = ~controlPi_13_1 & n616_ntk1;
  assign new_n2653_ = ~new_n2651_ & ~new_n2652_;
  assign new_n2654_ = ~controlPi_13_2 & new_n2653_;
  assign new_n2655_ = controlPi_13_1 & n673_ntk1;
  assign new_n2656_ = ~controlPi_13_1 & n664_ntk1;
  assign new_n2657_ = ~new_n2655_ & ~new_n2656_;
  assign new_n2658_ = controlPi_13_2 & new_n2657_;
  assign new_n2659_ = ~new_n2654_ & ~new_n2658_;
  assign new_n2660_ = controlPi_13_4 & ~new_n2659_;
  assign new_n2661_ = controlPi_13_1 & n457_ntk1;
  assign new_n2662_ = ~controlPi_13_1 & n454_ntk1;
  assign new_n2663_ = ~new_n2661_ & ~new_n2662_;
  assign new_n2664_ = ~controlPi_13_2 & new_n2663_;
  assign new_n2665_ = controlPi_13_1 & n507_ntk1;
  assign new_n2666_ = ~controlPi_13_1 & n468_ntk1;
  assign new_n2667_ = ~new_n2665_ & ~new_n2666_;
  assign new_n2668_ = controlPi_13_2 & new_n2667_;
  assign new_n2669_ = ~new_n2664_ & ~new_n2668_;
  assign new_n2670_ = ~controlPi_13_4 & ~new_n2669_;
  assign new_n2671_ = ~new_n2660_ & ~new_n2670_;
  assign new_n2672_ = ~controlPi_13_3 & ~new_n2671_;
  assign new_n2673_ = controlPi_13_1 & n600_ntk1;
  assign new_n2674_ = ~controlPi_13_1 & n582_ntk1;
  assign new_n2675_ = ~new_n2673_ & ~new_n2674_;
  assign new_n2676_ = controlPi_13_2 & new_n2675_;
  assign new_n2677_ = controlPi_13_1 & n525_ntk1;
  assign new_n2678_ = ~controlPi_13_1 & n511_ntk1;
  assign new_n2679_ = ~new_n2677_ & ~new_n2678_;
  assign new_n2680_ = ~controlPi_13_2 & new_n2679_;
  assign new_n2681_ = ~new_n2676_ & ~new_n2680_;
  assign new_n2682_ = controlPi_13_3 & ~new_n2681_;
  assign new_n2683_ = ~controlPi_13_4 & new_n2682_;
  assign new_n2684_ = ~new_n2672_ & ~new_n2683_;
  assign new_n2685_ = controlPi_13_5 & ~new_n2684_;
  assign new_n2686_ = ~new_n2650_ & ~new_n2685_;
  assign new_n2687_ = controlPi_13_0 & ~new_n2686_;
  assign new_n2688_ = ~controlPi_13_0 & new_n2686_;
  assign new_n2689_ = ~new_n2687_ & ~new_n2688_;
  assign new_n2690_ = ~new_n1946_ & ~new_n2689_;
  assign new_n2691_ = new_n1775_ & new_n2603_;
  assign new_n2692_ = new_n2690_ & ~new_n2691_;
  assign new_n2693_ = ~new_n2604_ & ~new_n2692_;
  assign new_n2694_ = ~controlPi_1_1 & ~n199_ntk1;
  assign new_n2695_ = controlPi_1_1 & ~n211_ntk1;
  assign new_n2696_ = ~new_n2694_ & ~new_n2695_;
  assign new_n2697_ = ~controlPi_1_2 & new_n2696_;
  assign new_n2698_ = ~controlPi_1_1 & ~n216_ntk1;
  assign new_n2699_ = controlPi_1_1 & ~n280_ntk1;
  assign new_n2700_ = ~new_n2698_ & ~new_n2699_;
  assign new_n2701_ = controlPi_1_2 & new_n2700_;
  assign new_n2702_ = ~new_n2697_ & ~new_n2701_;
  assign new_n2703_ = ~controlPi_1_3 & new_n2702_;
  assign new_n2704_ = ~controlPi_1_1 & ~n287_ntk1;
  assign new_n2705_ = controlPi_1_1 & ~n409_ntk1;
  assign new_n2706_ = ~new_n2704_ & ~new_n2705_;
  assign new_n2707_ = ~controlPi_1_2 & new_n2706_;
  assign new_n2708_ = ~controlPi_1_1 & ~n428_ntk1;
  assign new_n2709_ = controlPi_1_1 & ~n435_ntk1;
  assign new_n2710_ = ~new_n2708_ & ~new_n2709_;
  assign new_n2711_ = controlPi_1_2 & new_n2710_;
  assign new_n2712_ = ~new_n2707_ & ~new_n2711_;
  assign new_n2713_ = controlPi_1_3 & new_n2712_;
  assign new_n2714_ = ~new_n2703_ & ~new_n2713_;
  assign new_n2715_ = controlPi_1_4 & ~new_n2714_;
  assign new_n2716_ = ~controlPi_1_1 & ~n2_ntk1;
  assign new_n2717_ = controlPi_1_1 & ~n13_ntk1;
  assign new_n2718_ = ~new_n2716_ & ~new_n2717_;
  assign new_n2719_ = ~controlPi_1_2 & new_n2718_;
  assign new_n2720_ = ~controlPi_1_1 & ~n46_ntk1;
  assign new_n2721_ = controlPi_1_1 & ~n75_ntk1;
  assign new_n2722_ = ~new_n2720_ & ~new_n2721_;
  assign new_n2723_ = controlPi_1_2 & new_n2722_;
  assign new_n2724_ = ~new_n2719_ & ~new_n2723_;
  assign new_n2725_ = ~controlPi_1_3 & new_n2724_;
  assign new_n2726_ = ~controlPi_1_1 & ~n96_ntk1;
  assign new_n2727_ = controlPi_1_1 & ~n131_ntk1;
  assign new_n2728_ = ~new_n2726_ & ~new_n2727_;
  assign new_n2729_ = ~controlPi_1_2 & new_n2728_;
  assign new_n2730_ = ~controlPi_1_1 & ~n159_ntk1;
  assign new_n2731_ = controlPi_1_1 & ~n177_ntk1;
  assign new_n2732_ = ~new_n2730_ & ~new_n2731_;
  assign new_n2733_ = controlPi_1_2 & new_n2732_;
  assign new_n2734_ = ~new_n2729_ & ~new_n2733_;
  assign new_n2735_ = controlPi_1_3 & new_n2734_;
  assign new_n2736_ = ~new_n2725_ & ~new_n2735_;
  assign new_n2737_ = ~controlPi_1_4 & ~new_n2736_;
  assign new_n2738_ = ~new_n2715_ & ~new_n2737_;
  assign new_n2739_ = ~controlPi_1_5 & ~new_n2738_;
  assign new_n2740_ = controlPi_1_1 & n659_ntk1;
  assign new_n2741_ = ~controlPi_1_1 & n616_ntk1;
  assign new_n2742_ = ~new_n2740_ & ~new_n2741_;
  assign new_n2743_ = ~controlPi_1_2 & new_n2742_;
  assign new_n2744_ = controlPi_1_1 & n673_ntk1;
  assign new_n2745_ = ~controlPi_1_1 & n664_ntk1;
  assign new_n2746_ = ~new_n2744_ & ~new_n2745_;
  assign new_n2747_ = controlPi_1_2 & new_n2746_;
  assign new_n2748_ = ~new_n2743_ & ~new_n2747_;
  assign new_n2749_ = controlPi_1_4 & ~new_n2748_;
  assign new_n2750_ = controlPi_1_1 & n457_ntk1;
  assign new_n2751_ = ~controlPi_1_1 & n454_ntk1;
  assign new_n2752_ = ~new_n2750_ & ~new_n2751_;
  assign new_n2753_ = ~controlPi_1_2 & new_n2752_;
  assign new_n2754_ = controlPi_1_1 & n507_ntk1;
  assign new_n2755_ = ~controlPi_1_1 & n468_ntk1;
  assign new_n2756_ = ~new_n2754_ & ~new_n2755_;
  assign new_n2757_ = controlPi_1_2 & new_n2756_;
  assign new_n2758_ = ~new_n2753_ & ~new_n2757_;
  assign new_n2759_ = ~controlPi_1_4 & ~new_n2758_;
  assign new_n2760_ = ~new_n2749_ & ~new_n2759_;
  assign new_n2761_ = ~controlPi_1_3 & ~new_n2760_;
  assign new_n2762_ = controlPi_1_1 & n600_ntk1;
  assign new_n2763_ = ~controlPi_1_1 & n582_ntk1;
  assign new_n2764_ = ~new_n2762_ & ~new_n2763_;
  assign new_n2765_ = controlPi_1_2 & new_n2764_;
  assign new_n2766_ = controlPi_1_1 & n525_ntk1;
  assign new_n2767_ = ~controlPi_1_1 & n511_ntk1;
  assign new_n2768_ = ~new_n2766_ & ~new_n2767_;
  assign new_n2769_ = ~controlPi_1_2 & new_n2768_;
  assign new_n2770_ = ~new_n2765_ & ~new_n2769_;
  assign new_n2771_ = controlPi_1_3 & ~new_n2770_;
  assign new_n2772_ = ~controlPi_1_4 & new_n2771_;
  assign new_n2773_ = ~new_n2761_ & ~new_n2772_;
  assign new_n2774_ = controlPi_1_5 & ~new_n2773_;
  assign new_n2775_ = ~new_n2739_ & ~new_n2774_;
  assign new_n2776_ = controlPi_1_0 & ~new_n2775_;
  assign new_n2777_ = ~controlPi_1_0 & new_n2775_;
  assign new_n2778_ = ~new_n2776_ & ~new_n2777_;
  assign new_n2779_ = new_n2035_ & new_n2778_;
  assign new_n2780_ = ~new_n2035_ & ~new_n2778_;
  assign new_n2781_ = ~new_n2779_ & ~new_n2780_;
  assign new_n2782_ = new_n2693_ & ~new_n2781_;
  assign new_n2783_ = ~new_n2693_ & new_n2781_;
  assign new_n2784_ = ~new_n2782_ & ~new_n2783_;
  assign new_n2785_ = ~new_n2432_ & ~new_n2784_;
  assign new_n2786_ = ~new_n2518_ & ~new_n2785_;
  assign new_n2787_ = new_n2146_ & ~new_n2786_;
  assign new_n2788_ = ~new_n2413_ & ~new_n2787_;
  assign new_n2789_ = new_n1605_ & ~new_n2788_;
  assign new_n2790_ = ~new_n2127_ & ~new_n2789_;
  assign new_n2791_ = new_n1586_ & ~new_n2790_;
  assign new_n2792_ = ~new_n1110_ & ~new_n1281_;
  assign new_n2793_ = new_n1540_ & ~new_n2792_;
  assign new_n2794_ = ~new_n1540_ & new_n2792_;
  assign new_n2795_ = ~new_n2793_ & ~new_n2794_;
  assign new_n2796_ = ~new_n1586_ & ~new_n2795_;
  assign new_n2797_ = ~new_n2791_ & ~new_n2796_;
  assign new_n2798_ = new_n1567_ & ~new_n2797_;
  assign new_n2799_ = ~controlPi_41_1 & ~n199_ntk1;
  assign new_n2800_ = controlPi_41_1 & ~n211_ntk1;
  assign new_n2801_ = ~new_n2799_ & ~new_n2800_;
  assign new_n2802_ = ~controlPi_41_2 & new_n2801_;
  assign new_n2803_ = ~controlPi_41_1 & ~n216_ntk1;
  assign new_n2804_ = controlPi_41_1 & ~n280_ntk1;
  assign new_n2805_ = ~new_n2803_ & ~new_n2804_;
  assign new_n2806_ = controlPi_41_2 & new_n2805_;
  assign new_n2807_ = ~new_n2802_ & ~new_n2806_;
  assign new_n2808_ = ~controlPi_41_3 & new_n2807_;
  assign new_n2809_ = ~controlPi_41_1 & ~n287_ntk1;
  assign new_n2810_ = controlPi_41_1 & ~n409_ntk1;
  assign new_n2811_ = ~new_n2809_ & ~new_n2810_;
  assign new_n2812_ = ~controlPi_41_2 & new_n2811_;
  assign new_n2813_ = ~controlPi_41_1 & ~n428_ntk1;
  assign new_n2814_ = controlPi_41_1 & ~n435_ntk1;
  assign new_n2815_ = ~new_n2813_ & ~new_n2814_;
  assign new_n2816_ = controlPi_41_2 & new_n2815_;
  assign new_n2817_ = ~new_n2812_ & ~new_n2816_;
  assign new_n2818_ = controlPi_41_3 & new_n2817_;
  assign new_n2819_ = ~new_n2808_ & ~new_n2818_;
  assign new_n2820_ = controlPi_41_4 & ~new_n2819_;
  assign new_n2821_ = ~controlPi_41_1 & ~n2_ntk1;
  assign new_n2822_ = controlPi_41_1 & ~n13_ntk1;
  assign new_n2823_ = ~new_n2821_ & ~new_n2822_;
  assign new_n2824_ = ~controlPi_41_2 & new_n2823_;
  assign new_n2825_ = ~controlPi_41_1 & ~n46_ntk1;
  assign new_n2826_ = controlPi_41_1 & ~n75_ntk1;
  assign new_n2827_ = ~new_n2825_ & ~new_n2826_;
  assign new_n2828_ = controlPi_41_2 & new_n2827_;
  assign new_n2829_ = ~new_n2824_ & ~new_n2828_;
  assign new_n2830_ = ~controlPi_41_3 & new_n2829_;
  assign new_n2831_ = ~controlPi_41_1 & ~n96_ntk1;
  assign new_n2832_ = controlPi_41_1 & ~n131_ntk1;
  assign new_n2833_ = ~new_n2831_ & ~new_n2832_;
  assign new_n2834_ = ~controlPi_41_2 & new_n2833_;
  assign new_n2835_ = ~controlPi_41_1 & ~n159_ntk1;
  assign new_n2836_ = controlPi_41_1 & ~n177_ntk1;
  assign new_n2837_ = ~new_n2835_ & ~new_n2836_;
  assign new_n2838_ = controlPi_41_2 & new_n2837_;
  assign new_n2839_ = ~new_n2834_ & ~new_n2838_;
  assign new_n2840_ = controlPi_41_3 & new_n2839_;
  assign new_n2841_ = ~new_n2830_ & ~new_n2840_;
  assign new_n2842_ = ~controlPi_41_4 & ~new_n2841_;
  assign new_n2843_ = ~new_n2820_ & ~new_n2842_;
  assign new_n2844_ = ~controlPi_41_5 & ~new_n2843_;
  assign new_n2845_ = controlPi_41_1 & n659_ntk1;
  assign new_n2846_ = ~controlPi_41_1 & n616_ntk1;
  assign new_n2847_ = ~new_n2845_ & ~new_n2846_;
  assign new_n2848_ = ~controlPi_41_2 & new_n2847_;
  assign new_n2849_ = controlPi_41_1 & n673_ntk1;
  assign new_n2850_ = ~controlPi_41_1 & n664_ntk1;
  assign new_n2851_ = ~new_n2849_ & ~new_n2850_;
  assign new_n2852_ = controlPi_41_2 & new_n2851_;
  assign new_n2853_ = ~new_n2848_ & ~new_n2852_;
  assign new_n2854_ = controlPi_41_4 & ~new_n2853_;
  assign new_n2855_ = controlPi_41_1 & n457_ntk1;
  assign new_n2856_ = ~controlPi_41_1 & n454_ntk1;
  assign new_n2857_ = ~new_n2855_ & ~new_n2856_;
  assign new_n2858_ = ~controlPi_41_2 & new_n2857_;
  assign new_n2859_ = controlPi_41_1 & n507_ntk1;
  assign new_n2860_ = ~controlPi_41_1 & n468_ntk1;
  assign new_n2861_ = ~new_n2859_ & ~new_n2860_;
  assign new_n2862_ = controlPi_41_2 & new_n2861_;
  assign new_n2863_ = ~new_n2858_ & ~new_n2862_;
  assign new_n2864_ = ~controlPi_41_4 & ~new_n2863_;
  assign new_n2865_ = ~new_n2854_ & ~new_n2864_;
  assign new_n2866_ = ~controlPi_41_3 & ~new_n2865_;
  assign new_n2867_ = controlPi_41_1 & n600_ntk1;
  assign new_n2868_ = ~controlPi_41_1 & n582_ntk1;
  assign new_n2869_ = ~new_n2867_ & ~new_n2868_;
  assign new_n2870_ = controlPi_41_2 & new_n2869_;
  assign new_n2871_ = controlPi_41_1 & n525_ntk1;
  assign new_n2872_ = ~controlPi_41_1 & n511_ntk1;
  assign new_n2873_ = ~new_n2871_ & ~new_n2872_;
  assign new_n2874_ = ~controlPi_41_2 & new_n2873_;
  assign new_n2875_ = ~new_n2870_ & ~new_n2874_;
  assign new_n2876_ = controlPi_41_3 & ~new_n2875_;
  assign new_n2877_ = ~controlPi_41_4 & new_n2876_;
  assign new_n2878_ = ~new_n2866_ & ~new_n2877_;
  assign new_n2879_ = controlPi_41_5 & ~new_n2878_;
  assign new_n2880_ = ~new_n2844_ & ~new_n2879_;
  assign new_n2881_ = controlPi_41_0 & ~new_n2880_;
  assign new_n2882_ = ~controlPi_41_0 & new_n2880_;
  assign new_n2883_ = ~new_n2881_ & ~new_n2882_;
  assign new_n2884_ = ~controlPi_25_1 & ~n199_ntk1;
  assign new_n2885_ = controlPi_25_1 & ~n211_ntk1;
  assign new_n2886_ = ~new_n2884_ & ~new_n2885_;
  assign new_n2887_ = ~controlPi_25_2 & new_n2886_;
  assign new_n2888_ = ~controlPi_25_1 & ~n216_ntk1;
  assign new_n2889_ = controlPi_25_1 & ~n280_ntk1;
  assign new_n2890_ = ~new_n2888_ & ~new_n2889_;
  assign new_n2891_ = controlPi_25_2 & new_n2890_;
  assign new_n2892_ = ~new_n2887_ & ~new_n2891_;
  assign new_n2893_ = ~controlPi_25_3 & new_n2892_;
  assign new_n2894_ = ~controlPi_25_1 & ~n287_ntk1;
  assign new_n2895_ = controlPi_25_1 & ~n409_ntk1;
  assign new_n2896_ = ~new_n2894_ & ~new_n2895_;
  assign new_n2897_ = ~controlPi_25_2 & new_n2896_;
  assign new_n2898_ = ~controlPi_25_1 & ~n428_ntk1;
  assign new_n2899_ = controlPi_25_1 & ~n435_ntk1;
  assign new_n2900_ = ~new_n2898_ & ~new_n2899_;
  assign new_n2901_ = controlPi_25_2 & new_n2900_;
  assign new_n2902_ = ~new_n2897_ & ~new_n2901_;
  assign new_n2903_ = controlPi_25_3 & new_n2902_;
  assign new_n2904_ = ~new_n2893_ & ~new_n2903_;
  assign new_n2905_ = controlPi_25_4 & ~new_n2904_;
  assign new_n2906_ = ~controlPi_25_1 & ~n2_ntk1;
  assign new_n2907_ = controlPi_25_1 & ~n13_ntk1;
  assign new_n2908_ = ~new_n2906_ & ~new_n2907_;
  assign new_n2909_ = ~controlPi_25_2 & new_n2908_;
  assign new_n2910_ = ~controlPi_25_1 & ~n46_ntk1;
  assign new_n2911_ = controlPi_25_1 & ~n75_ntk1;
  assign new_n2912_ = ~new_n2910_ & ~new_n2911_;
  assign new_n2913_ = controlPi_25_2 & new_n2912_;
  assign new_n2914_ = ~new_n2909_ & ~new_n2913_;
  assign new_n2915_ = ~controlPi_25_3 & new_n2914_;
  assign new_n2916_ = ~controlPi_25_1 & ~n96_ntk1;
  assign new_n2917_ = controlPi_25_1 & ~n131_ntk1;
  assign new_n2918_ = ~new_n2916_ & ~new_n2917_;
  assign new_n2919_ = ~controlPi_25_2 & new_n2918_;
  assign new_n2920_ = ~controlPi_25_1 & ~n159_ntk1;
  assign new_n2921_ = controlPi_25_1 & ~n177_ntk1;
  assign new_n2922_ = ~new_n2920_ & ~new_n2921_;
  assign new_n2923_ = controlPi_25_2 & new_n2922_;
  assign new_n2924_ = ~new_n2919_ & ~new_n2923_;
  assign new_n2925_ = controlPi_25_3 & new_n2924_;
  assign new_n2926_ = ~new_n2915_ & ~new_n2925_;
  assign new_n2927_ = ~controlPi_25_4 & ~new_n2926_;
  assign new_n2928_ = ~new_n2905_ & ~new_n2927_;
  assign new_n2929_ = ~controlPi_25_5 & ~new_n2928_;
  assign new_n2930_ = controlPi_25_1 & n659_ntk1;
  assign new_n2931_ = ~controlPi_25_1 & n616_ntk1;
  assign new_n2932_ = ~new_n2930_ & ~new_n2931_;
  assign new_n2933_ = ~controlPi_25_2 & new_n2932_;
  assign new_n2934_ = controlPi_25_1 & n673_ntk1;
  assign new_n2935_ = ~controlPi_25_1 & n664_ntk1;
  assign new_n2936_ = ~new_n2934_ & ~new_n2935_;
  assign new_n2937_ = controlPi_25_2 & new_n2936_;
  assign new_n2938_ = ~new_n2933_ & ~new_n2937_;
  assign new_n2939_ = controlPi_25_4 & ~new_n2938_;
  assign new_n2940_ = controlPi_25_1 & n457_ntk1;
  assign new_n2941_ = ~controlPi_25_1 & n454_ntk1;
  assign new_n2942_ = ~new_n2940_ & ~new_n2941_;
  assign new_n2943_ = ~controlPi_25_2 & new_n2942_;
  assign new_n2944_ = controlPi_25_1 & n507_ntk1;
  assign new_n2945_ = ~controlPi_25_1 & n468_ntk1;
  assign new_n2946_ = ~new_n2944_ & ~new_n2945_;
  assign new_n2947_ = controlPi_25_2 & new_n2946_;
  assign new_n2948_ = ~new_n2943_ & ~new_n2947_;
  assign new_n2949_ = ~controlPi_25_4 & ~new_n2948_;
  assign new_n2950_ = ~new_n2939_ & ~new_n2949_;
  assign new_n2951_ = ~controlPi_25_3 & ~new_n2950_;
  assign new_n2952_ = controlPi_25_1 & n600_ntk1;
  assign new_n2953_ = ~controlPi_25_1 & n582_ntk1;
  assign new_n2954_ = ~new_n2952_ & ~new_n2953_;
  assign new_n2955_ = controlPi_25_2 & new_n2954_;
  assign new_n2956_ = controlPi_25_1 & n525_ntk1;
  assign new_n2957_ = ~controlPi_25_1 & n511_ntk1;
  assign new_n2958_ = ~new_n2956_ & ~new_n2957_;
  assign new_n2959_ = ~controlPi_25_2 & new_n2958_;
  assign new_n2960_ = ~new_n2955_ & ~new_n2959_;
  assign new_n2961_ = controlPi_25_3 & ~new_n2960_;
  assign new_n2962_ = ~controlPi_25_4 & new_n2961_;
  assign new_n2963_ = ~new_n2951_ & ~new_n2962_;
  assign new_n2964_ = controlPi_25_5 & ~new_n2963_;
  assign new_n2965_ = ~new_n2929_ & ~new_n2964_;
  assign new_n2966_ = controlPi_25_0 & ~new_n2965_;
  assign new_n2967_ = ~controlPi_25_0 & new_n2965_;
  assign new_n2968_ = ~new_n2966_ & ~new_n2967_;
  assign new_n2969_ = ~new_n2883_ & new_n2968_;
  assign new_n2970_ = new_n2883_ & ~new_n2968_;
  assign new_n2971_ = ~new_n2969_ & ~new_n2970_;
  assign new_n2972_ = ~new_n1110_ & ~new_n2883_;
  assign new_n2973_ = ~new_n1540_ & new_n2972_;
  assign new_n2974_ = new_n1540_ & ~new_n2972_;
  assign new_n2975_ = ~new_n2973_ & ~new_n2974_;
  assign new_n2976_ = ~new_n2971_ & ~new_n2975_;
  assign new_n2977_ = new_n2971_ & new_n2975_;
  assign new_n2978_ = ~new_n2976_ & ~new_n2977_;
  assign new_n2979_ = ~new_n1567_ & new_n2978_;
  assign new_n2980_ = ~new_n2798_ & ~new_n2979_;
  assign new_n2981_ = ~new_n1548_ & ~new_n2980_;
  assign new_n2982_ = new_n1548_ & new_n2980_;
  assign new_n2983_ = ~new_n2981_ & ~new_n2982_;
  assign new_n2984_ = ~controlPi_63_1 & ~n199_ntk1;
  assign new_n2985_ = controlPi_63_1 & ~n211_ntk1;
  assign new_n2986_ = ~new_n2984_ & ~new_n2985_;
  assign new_n2987_ = ~controlPi_63_2 & new_n2986_;
  assign new_n2988_ = ~controlPi_63_1 & ~n216_ntk1;
  assign new_n2989_ = controlPi_63_1 & ~n280_ntk1;
  assign new_n2990_ = ~new_n2988_ & ~new_n2989_;
  assign new_n2991_ = controlPi_63_2 & new_n2990_;
  assign new_n2992_ = ~new_n2987_ & ~new_n2991_;
  assign new_n2993_ = ~controlPi_63_3 & new_n2992_;
  assign new_n2994_ = ~controlPi_63_1 & ~n287_ntk1;
  assign new_n2995_ = controlPi_63_1 & ~n409_ntk1;
  assign new_n2996_ = ~new_n2994_ & ~new_n2995_;
  assign new_n2997_ = ~controlPi_63_2 & new_n2996_;
  assign new_n2998_ = ~controlPi_63_1 & ~n428_ntk1;
  assign new_n2999_ = controlPi_63_1 & ~n435_ntk1;
  assign new_n3000_ = ~new_n2998_ & ~new_n2999_;
  assign new_n3001_ = controlPi_63_2 & new_n3000_;
  assign new_n3002_ = ~new_n2997_ & ~new_n3001_;
  assign new_n3003_ = controlPi_63_3 & new_n3002_;
  assign new_n3004_ = ~new_n2993_ & ~new_n3003_;
  assign new_n3005_ = controlPi_63_4 & ~new_n3004_;
  assign new_n3006_ = ~controlPi_63_1 & ~n2_ntk1;
  assign new_n3007_ = controlPi_63_1 & ~n13_ntk1;
  assign new_n3008_ = ~new_n3006_ & ~new_n3007_;
  assign new_n3009_ = ~controlPi_63_2 & new_n3008_;
  assign new_n3010_ = ~controlPi_63_1 & ~n46_ntk1;
  assign new_n3011_ = controlPi_63_1 & ~n75_ntk1;
  assign new_n3012_ = ~new_n3010_ & ~new_n3011_;
  assign new_n3013_ = controlPi_63_2 & new_n3012_;
  assign new_n3014_ = ~new_n3009_ & ~new_n3013_;
  assign new_n3015_ = ~controlPi_63_3 & new_n3014_;
  assign new_n3016_ = ~controlPi_63_1 & ~n96_ntk1;
  assign new_n3017_ = controlPi_63_1 & ~n131_ntk1;
  assign new_n3018_ = ~new_n3016_ & ~new_n3017_;
  assign new_n3019_ = ~controlPi_63_2 & new_n3018_;
  assign new_n3020_ = ~controlPi_63_1 & ~n159_ntk1;
  assign new_n3021_ = controlPi_63_1 & ~n177_ntk1;
  assign new_n3022_ = ~new_n3020_ & ~new_n3021_;
  assign new_n3023_ = controlPi_63_2 & new_n3022_;
  assign new_n3024_ = ~new_n3019_ & ~new_n3023_;
  assign new_n3025_ = controlPi_63_3 & new_n3024_;
  assign new_n3026_ = ~new_n3015_ & ~new_n3025_;
  assign new_n3027_ = ~controlPi_63_4 & ~new_n3026_;
  assign new_n3028_ = ~new_n3005_ & ~new_n3027_;
  assign new_n3029_ = ~controlPi_63_5 & ~new_n3028_;
  assign new_n3030_ = controlPi_63_1 & n659_ntk1;
  assign new_n3031_ = ~controlPi_63_1 & n616_ntk1;
  assign new_n3032_ = ~new_n3030_ & ~new_n3031_;
  assign new_n3033_ = ~controlPi_63_2 & new_n3032_;
  assign new_n3034_ = controlPi_63_1 & n673_ntk1;
  assign new_n3035_ = ~controlPi_63_1 & n664_ntk1;
  assign new_n3036_ = ~new_n3034_ & ~new_n3035_;
  assign new_n3037_ = controlPi_63_2 & new_n3036_;
  assign new_n3038_ = ~new_n3033_ & ~new_n3037_;
  assign new_n3039_ = controlPi_63_4 & ~new_n3038_;
  assign new_n3040_ = controlPi_63_1 & n457_ntk1;
  assign new_n3041_ = ~controlPi_63_1 & n454_ntk1;
  assign new_n3042_ = ~new_n3040_ & ~new_n3041_;
  assign new_n3043_ = ~controlPi_63_2 & new_n3042_;
  assign new_n3044_ = controlPi_63_1 & n507_ntk1;
  assign new_n3045_ = ~controlPi_63_1 & n468_ntk1;
  assign new_n3046_ = ~new_n3044_ & ~new_n3045_;
  assign new_n3047_ = controlPi_63_2 & new_n3046_;
  assign new_n3048_ = ~new_n3043_ & ~new_n3047_;
  assign new_n3049_ = ~controlPi_63_4 & ~new_n3048_;
  assign new_n3050_ = ~new_n3039_ & ~new_n3049_;
  assign new_n3051_ = ~controlPi_63_3 & ~new_n3050_;
  assign new_n3052_ = controlPi_63_1 & n600_ntk1;
  assign new_n3053_ = ~controlPi_63_1 & n582_ntk1;
  assign new_n3054_ = ~new_n3052_ & ~new_n3053_;
  assign new_n3055_ = controlPi_63_2 & new_n3054_;
  assign new_n3056_ = controlPi_63_1 & n525_ntk1;
  assign new_n3057_ = ~controlPi_63_1 & n511_ntk1;
  assign new_n3058_ = ~new_n3056_ & ~new_n3057_;
  assign new_n3059_ = ~controlPi_63_2 & new_n3058_;
  assign new_n3060_ = ~new_n3055_ & ~new_n3059_;
  assign new_n3061_ = controlPi_63_3 & ~new_n3060_;
  assign new_n3062_ = ~controlPi_63_4 & new_n3061_;
  assign new_n3063_ = ~new_n3051_ & ~new_n3062_;
  assign new_n3064_ = controlPi_63_5 & ~new_n3063_;
  assign new_n3065_ = ~new_n3029_ & ~new_n3064_;
  assign new_n3066_ = controlPi_63_0 & ~new_n3065_;
  assign new_n3067_ = ~controlPi_63_0 & new_n3065_;
  assign new_n3068_ = ~new_n3066_ & ~new_n3067_;
  assign new_n3069_ = new_n939_ & ~new_n3068_;
  assign new_n3070_ = ~new_n1196_ & ~new_n1368_;
  assign new_n3071_ = new_n1367_ & ~new_n3070_;
  assign new_n3072_ = ~new_n1367_ & new_n3070_;
  assign new_n3073_ = ~new_n3071_ & ~new_n3072_;
  assign new_n3074_ = ~new_n939_ & ~new_n3073_;
  assign new_n3075_ = ~new_n3069_ & ~new_n3074_;
  assign new_n3076_ = new_n1110_ & new_n2883_;
  assign new_n3077_ = ~new_n2972_ & ~new_n3076_;
  assign new_n3078_ = ~new_n1567_ & new_n3077_;
  assign new_n3079_ = new_n1110_ & new_n1281_;
  assign new_n3080_ = ~new_n1586_ & ~new_n3079_;
  assign new_n3081_ = ~new_n2792_ & new_n3080_;
  assign new_n3082_ = ~controlPi_56_1 & ~n199_ntk1;
  assign new_n3083_ = controlPi_56_1 & ~n211_ntk1;
  assign new_n3084_ = ~new_n3082_ & ~new_n3083_;
  assign new_n3085_ = ~controlPi_56_2 & new_n3084_;
  assign new_n3086_ = ~controlPi_56_1 & ~n216_ntk1;
  assign new_n3087_ = controlPi_56_1 & ~n280_ntk1;
  assign new_n3088_ = ~new_n3086_ & ~new_n3087_;
  assign new_n3089_ = controlPi_56_2 & new_n3088_;
  assign new_n3090_ = ~new_n3085_ & ~new_n3089_;
  assign new_n3091_ = ~controlPi_56_3 & new_n3090_;
  assign new_n3092_ = ~controlPi_56_1 & ~n287_ntk1;
  assign new_n3093_ = controlPi_56_1 & ~n409_ntk1;
  assign new_n3094_ = ~new_n3092_ & ~new_n3093_;
  assign new_n3095_ = ~controlPi_56_2 & new_n3094_;
  assign new_n3096_ = ~controlPi_56_1 & ~n428_ntk1;
  assign new_n3097_ = controlPi_56_1 & ~n435_ntk1;
  assign new_n3098_ = ~new_n3096_ & ~new_n3097_;
  assign new_n3099_ = controlPi_56_2 & new_n3098_;
  assign new_n3100_ = ~new_n3095_ & ~new_n3099_;
  assign new_n3101_ = controlPi_56_3 & new_n3100_;
  assign new_n3102_ = ~new_n3091_ & ~new_n3101_;
  assign new_n3103_ = controlPi_56_4 & ~new_n3102_;
  assign new_n3104_ = ~controlPi_56_1 & ~n2_ntk1;
  assign new_n3105_ = controlPi_56_1 & ~n13_ntk1;
  assign new_n3106_ = ~new_n3104_ & ~new_n3105_;
  assign new_n3107_ = ~controlPi_56_2 & new_n3106_;
  assign new_n3108_ = ~controlPi_56_1 & ~n46_ntk1;
  assign new_n3109_ = controlPi_56_1 & ~n75_ntk1;
  assign new_n3110_ = ~new_n3108_ & ~new_n3109_;
  assign new_n3111_ = controlPi_56_2 & new_n3110_;
  assign new_n3112_ = ~new_n3107_ & ~new_n3111_;
  assign new_n3113_ = ~controlPi_56_3 & new_n3112_;
  assign new_n3114_ = ~controlPi_56_1 & ~n96_ntk1;
  assign new_n3115_ = controlPi_56_1 & ~n131_ntk1;
  assign new_n3116_ = ~new_n3114_ & ~new_n3115_;
  assign new_n3117_ = ~controlPi_56_2 & new_n3116_;
  assign new_n3118_ = ~controlPi_56_1 & ~n159_ntk1;
  assign new_n3119_ = controlPi_56_1 & ~n177_ntk1;
  assign new_n3120_ = ~new_n3118_ & ~new_n3119_;
  assign new_n3121_ = controlPi_56_2 & new_n3120_;
  assign new_n3122_ = ~new_n3117_ & ~new_n3121_;
  assign new_n3123_ = controlPi_56_3 & new_n3122_;
  assign new_n3124_ = ~new_n3113_ & ~new_n3123_;
  assign new_n3125_ = ~controlPi_56_4 & ~new_n3124_;
  assign new_n3126_ = ~new_n3103_ & ~new_n3125_;
  assign new_n3127_ = ~controlPi_56_5 & ~new_n3126_;
  assign new_n3128_ = controlPi_56_1 & n659_ntk1;
  assign new_n3129_ = ~controlPi_56_1 & n616_ntk1;
  assign new_n3130_ = ~new_n3128_ & ~new_n3129_;
  assign new_n3131_ = ~controlPi_56_2 & new_n3130_;
  assign new_n3132_ = controlPi_56_1 & n673_ntk1;
  assign new_n3133_ = ~controlPi_56_1 & n664_ntk1;
  assign new_n3134_ = ~new_n3132_ & ~new_n3133_;
  assign new_n3135_ = controlPi_56_2 & new_n3134_;
  assign new_n3136_ = ~new_n3131_ & ~new_n3135_;
  assign new_n3137_ = controlPi_56_4 & ~new_n3136_;
  assign new_n3138_ = controlPi_56_1 & n457_ntk1;
  assign new_n3139_ = ~controlPi_56_1 & n454_ntk1;
  assign new_n3140_ = ~new_n3138_ & ~new_n3139_;
  assign new_n3141_ = ~controlPi_56_2 & new_n3140_;
  assign new_n3142_ = controlPi_56_1 & n507_ntk1;
  assign new_n3143_ = ~controlPi_56_1 & n468_ntk1;
  assign new_n3144_ = ~new_n3142_ & ~new_n3143_;
  assign new_n3145_ = controlPi_56_2 & new_n3144_;
  assign new_n3146_ = ~new_n3141_ & ~new_n3145_;
  assign new_n3147_ = ~controlPi_56_4 & ~new_n3146_;
  assign new_n3148_ = ~new_n3137_ & ~new_n3147_;
  assign new_n3149_ = ~controlPi_56_3 & ~new_n3148_;
  assign new_n3150_ = controlPi_56_1 & n600_ntk1;
  assign new_n3151_ = ~controlPi_56_1 & n582_ntk1;
  assign new_n3152_ = ~new_n3150_ & ~new_n3151_;
  assign new_n3153_ = controlPi_56_2 & new_n3152_;
  assign new_n3154_ = controlPi_56_1 & n525_ntk1;
  assign new_n3155_ = ~controlPi_56_1 & n511_ntk1;
  assign new_n3156_ = ~new_n3154_ & ~new_n3155_;
  assign new_n3157_ = ~controlPi_56_2 & new_n3156_;
  assign new_n3158_ = ~new_n3153_ & ~new_n3157_;
  assign new_n3159_ = controlPi_56_3 & ~new_n3158_;
  assign new_n3160_ = ~controlPi_56_4 & new_n3159_;
  assign new_n3161_ = ~new_n3149_ & ~new_n3160_;
  assign new_n3162_ = controlPi_56_5 & ~new_n3161_;
  assign new_n3163_ = ~new_n3127_ & ~new_n3162_;
  assign new_n3164_ = controlPi_56_0 & ~new_n3163_;
  assign new_n3165_ = ~controlPi_56_0 & new_n3163_;
  assign new_n3166_ = ~new_n3164_ & ~new_n3165_;
  assign new_n3167_ = new_n2432_ & ~new_n3166_;
  assign new_n3168_ = ~new_n2604_ & ~new_n2691_;
  assign new_n3169_ = new_n2690_ & ~new_n3168_;
  assign new_n3170_ = ~new_n2690_ & new_n3168_;
  assign new_n3171_ = ~new_n3169_ & ~new_n3170_;
  assign new_n3172_ = ~new_n2432_ & ~new_n3171_;
  assign new_n3173_ = ~new_n3167_ & ~new_n3172_;
  assign new_n3174_ = new_n2146_ & new_n3173_;
  assign new_n3175_ = ~new_n2232_ & ~new_n2319_;
  assign new_n3176_ = new_n2318_ & ~new_n3175_;
  assign new_n3177_ = ~new_n2318_ & new_n3175_;
  assign new_n3178_ = ~new_n3176_ & ~new_n3177_;
  assign new_n3179_ = ~new_n2146_ & new_n3178_;
  assign new_n3180_ = ~new_n3174_ & ~new_n3179_;
  assign new_n3181_ = new_n1605_ & ~new_n3180_;
  assign new_n3182_ = ~new_n1776_ & ~new_n1948_;
  assign new_n3183_ = new_n1947_ & ~new_n3182_;
  assign new_n3184_ = ~new_n1947_ & new_n3182_;
  assign new_n3185_ = ~new_n3183_ & ~new_n3184_;
  assign new_n3186_ = ~new_n1605_ & new_n3185_;
  assign new_n3187_ = new_n1586_ & ~new_n3186_;
  assign new_n3188_ = ~new_n3181_ & new_n3187_;
  assign new_n3189_ = ~new_n3081_ & ~new_n3188_;
  assign new_n3190_ = new_n1567_ & ~new_n3189_;
  assign new_n3191_ = ~new_n3078_ & ~new_n3190_;
  assign new_n3192_ = ~controlPi_72_1 & ~n199_ntk1;
  assign new_n3193_ = controlPi_72_1 & ~n211_ntk1;
  assign new_n3194_ = ~new_n3192_ & ~new_n3193_;
  assign new_n3195_ = ~controlPi_72_2 & new_n3194_;
  assign new_n3196_ = ~controlPi_72_1 & ~n216_ntk1;
  assign new_n3197_ = controlPi_72_1 & ~n280_ntk1;
  assign new_n3198_ = ~new_n3196_ & ~new_n3197_;
  assign new_n3199_ = controlPi_72_2 & new_n3198_;
  assign new_n3200_ = ~new_n3195_ & ~new_n3199_;
  assign new_n3201_ = ~controlPi_72_3 & new_n3200_;
  assign new_n3202_ = ~controlPi_72_1 & ~n287_ntk1;
  assign new_n3203_ = controlPi_72_1 & ~n409_ntk1;
  assign new_n3204_ = ~new_n3202_ & ~new_n3203_;
  assign new_n3205_ = ~controlPi_72_2 & new_n3204_;
  assign new_n3206_ = ~controlPi_72_1 & ~n428_ntk1;
  assign new_n3207_ = controlPi_72_1 & ~n435_ntk1;
  assign new_n3208_ = ~new_n3206_ & ~new_n3207_;
  assign new_n3209_ = controlPi_72_2 & new_n3208_;
  assign new_n3210_ = ~new_n3205_ & ~new_n3209_;
  assign new_n3211_ = controlPi_72_3 & new_n3210_;
  assign new_n3212_ = ~new_n3201_ & ~new_n3211_;
  assign new_n3213_ = controlPi_72_4 & ~new_n3212_;
  assign new_n3214_ = ~controlPi_72_1 & ~n2_ntk1;
  assign new_n3215_ = controlPi_72_1 & ~n13_ntk1;
  assign new_n3216_ = ~new_n3214_ & ~new_n3215_;
  assign new_n3217_ = ~controlPi_72_2 & new_n3216_;
  assign new_n3218_ = ~controlPi_72_1 & ~n46_ntk1;
  assign new_n3219_ = controlPi_72_1 & ~n75_ntk1;
  assign new_n3220_ = ~new_n3218_ & ~new_n3219_;
  assign new_n3221_ = controlPi_72_2 & new_n3220_;
  assign new_n3222_ = ~new_n3217_ & ~new_n3221_;
  assign new_n3223_ = ~controlPi_72_3 & new_n3222_;
  assign new_n3224_ = ~controlPi_72_1 & ~n96_ntk1;
  assign new_n3225_ = controlPi_72_1 & ~n131_ntk1;
  assign new_n3226_ = ~new_n3224_ & ~new_n3225_;
  assign new_n3227_ = ~controlPi_72_2 & new_n3226_;
  assign new_n3228_ = ~controlPi_72_1 & ~n159_ntk1;
  assign new_n3229_ = controlPi_72_1 & ~n177_ntk1;
  assign new_n3230_ = ~new_n3228_ & ~new_n3229_;
  assign new_n3231_ = controlPi_72_2 & new_n3230_;
  assign new_n3232_ = ~new_n3227_ & ~new_n3231_;
  assign new_n3233_ = controlPi_72_3 & new_n3232_;
  assign new_n3234_ = ~new_n3223_ & ~new_n3233_;
  assign new_n3235_ = ~controlPi_72_4 & ~new_n3234_;
  assign new_n3236_ = ~new_n3213_ & ~new_n3235_;
  assign new_n3237_ = ~controlPi_72_5 & ~new_n3236_;
  assign new_n3238_ = controlPi_72_1 & n659_ntk1;
  assign new_n3239_ = ~controlPi_72_1 & n616_ntk1;
  assign new_n3240_ = ~new_n3238_ & ~new_n3239_;
  assign new_n3241_ = ~controlPi_72_2 & new_n3240_;
  assign new_n3242_ = controlPi_72_1 & n673_ntk1;
  assign new_n3243_ = ~controlPi_72_1 & n664_ntk1;
  assign new_n3244_ = ~new_n3242_ & ~new_n3243_;
  assign new_n3245_ = controlPi_72_2 & new_n3244_;
  assign new_n3246_ = ~new_n3241_ & ~new_n3245_;
  assign new_n3247_ = controlPi_72_4 & ~new_n3246_;
  assign new_n3248_ = controlPi_72_1 & n457_ntk1;
  assign new_n3249_ = ~controlPi_72_1 & n454_ntk1;
  assign new_n3250_ = ~new_n3248_ & ~new_n3249_;
  assign new_n3251_ = ~controlPi_72_2 & new_n3250_;
  assign new_n3252_ = controlPi_72_1 & n507_ntk1;
  assign new_n3253_ = ~controlPi_72_1 & n468_ntk1;
  assign new_n3254_ = ~new_n3252_ & ~new_n3253_;
  assign new_n3255_ = controlPi_72_2 & new_n3254_;
  assign new_n3256_ = ~new_n3251_ & ~new_n3255_;
  assign new_n3257_ = ~controlPi_72_4 & ~new_n3256_;
  assign new_n3258_ = ~new_n3247_ & ~new_n3257_;
  assign new_n3259_ = ~controlPi_72_3 & ~new_n3258_;
  assign new_n3260_ = controlPi_72_1 & n600_ntk1;
  assign new_n3261_ = ~controlPi_72_1 & n582_ntk1;
  assign new_n3262_ = ~new_n3260_ & ~new_n3261_;
  assign new_n3263_ = controlPi_72_2 & new_n3262_;
  assign new_n3264_ = controlPi_72_1 & n525_ntk1;
  assign new_n3265_ = ~controlPi_72_1 & n511_ntk1;
  assign new_n3266_ = ~new_n3264_ & ~new_n3265_;
  assign new_n3267_ = ~controlPi_72_2 & new_n3266_;
  assign new_n3268_ = ~new_n3263_ & ~new_n3267_;
  assign new_n3269_ = controlPi_72_3 & ~new_n3268_;
  assign new_n3270_ = ~controlPi_72_4 & new_n3269_;
  assign new_n3271_ = ~new_n3259_ & ~new_n3270_;
  assign new_n3272_ = controlPi_72_5 & ~new_n3271_;
  assign new_n3273_ = ~new_n3237_ & ~new_n3272_;
  assign new_n3274_ = controlPi_72_0 & ~new_n3273_;
  assign new_n3275_ = ~controlPi_72_0 & new_n3273_;
  assign new_n3276_ = ~new_n3274_ & ~new_n3275_;
  assign new_n3277_ = new_n939_ & ~new_n3276_;
  assign new_n3278_ = new_n1281_ & new_n1366_;
  assign new_n3279_ = ~new_n1367_ & ~new_n3278_;
  assign new_n3280_ = ~new_n939_ & new_n3279_;
  assign new_n3281_ = ~new_n3277_ & ~new_n3280_;
  assign new_n3282_ = ~new_n1281_ & ~new_n1586_;
  assign new_n3283_ = new_n1861_ & new_n1946_;
  assign new_n3284_ = ~new_n1947_ & ~new_n3283_;
  assign new_n3285_ = ~new_n1605_ & ~new_n3284_;
  assign new_n3286_ = ~controlPi_35_1 & ~n199_ntk1;
  assign new_n3287_ = controlPi_35_1 & ~n211_ntk1;
  assign new_n3288_ = ~new_n3286_ & ~new_n3287_;
  assign new_n3289_ = ~controlPi_35_2 & new_n3288_;
  assign new_n3290_ = ~controlPi_35_1 & ~n216_ntk1;
  assign new_n3291_ = controlPi_35_1 & ~n280_ntk1;
  assign new_n3292_ = ~new_n3290_ & ~new_n3291_;
  assign new_n3293_ = controlPi_35_2 & new_n3292_;
  assign new_n3294_ = ~new_n3289_ & ~new_n3293_;
  assign new_n3295_ = ~controlPi_35_3 & new_n3294_;
  assign new_n3296_ = ~controlPi_35_1 & ~n287_ntk1;
  assign new_n3297_ = controlPi_35_1 & ~n409_ntk1;
  assign new_n3298_ = ~new_n3296_ & ~new_n3297_;
  assign new_n3299_ = ~controlPi_35_2 & new_n3298_;
  assign new_n3300_ = ~controlPi_35_1 & ~n428_ntk1;
  assign new_n3301_ = controlPi_35_1 & ~n435_ntk1;
  assign new_n3302_ = ~new_n3300_ & ~new_n3301_;
  assign new_n3303_ = controlPi_35_2 & new_n3302_;
  assign new_n3304_ = ~new_n3299_ & ~new_n3303_;
  assign new_n3305_ = controlPi_35_3 & new_n3304_;
  assign new_n3306_ = ~new_n3295_ & ~new_n3305_;
  assign new_n3307_ = controlPi_35_4 & ~new_n3306_;
  assign new_n3308_ = ~controlPi_35_1 & ~n2_ntk1;
  assign new_n3309_ = controlPi_35_1 & ~n13_ntk1;
  assign new_n3310_ = ~new_n3308_ & ~new_n3309_;
  assign new_n3311_ = ~controlPi_35_2 & new_n3310_;
  assign new_n3312_ = ~controlPi_35_1 & ~n46_ntk1;
  assign new_n3313_ = controlPi_35_1 & ~n75_ntk1;
  assign new_n3314_ = ~new_n3312_ & ~new_n3313_;
  assign new_n3315_ = controlPi_35_2 & new_n3314_;
  assign new_n3316_ = ~new_n3311_ & ~new_n3315_;
  assign new_n3317_ = ~controlPi_35_3 & new_n3316_;
  assign new_n3318_ = ~controlPi_35_1 & ~n96_ntk1;
  assign new_n3319_ = controlPi_35_1 & ~n131_ntk1;
  assign new_n3320_ = ~new_n3318_ & ~new_n3319_;
  assign new_n3321_ = ~controlPi_35_2 & new_n3320_;
  assign new_n3322_ = ~controlPi_35_1 & ~n159_ntk1;
  assign new_n3323_ = controlPi_35_1 & ~n177_ntk1;
  assign new_n3324_ = ~new_n3322_ & ~new_n3323_;
  assign new_n3325_ = controlPi_35_2 & new_n3324_;
  assign new_n3326_ = ~new_n3321_ & ~new_n3325_;
  assign new_n3327_ = controlPi_35_3 & new_n3326_;
  assign new_n3328_ = ~new_n3317_ & ~new_n3327_;
  assign new_n3329_ = ~controlPi_35_4 & ~new_n3328_;
  assign new_n3330_ = ~new_n3307_ & ~new_n3329_;
  assign new_n3331_ = ~controlPi_35_5 & ~new_n3330_;
  assign new_n3332_ = controlPi_35_1 & n659_ntk1;
  assign new_n3333_ = ~controlPi_35_1 & n616_ntk1;
  assign new_n3334_ = ~new_n3332_ & ~new_n3333_;
  assign new_n3335_ = ~controlPi_35_2 & new_n3334_;
  assign new_n3336_ = controlPi_35_1 & n673_ntk1;
  assign new_n3337_ = ~controlPi_35_1 & n664_ntk1;
  assign new_n3338_ = ~new_n3336_ & ~new_n3337_;
  assign new_n3339_ = controlPi_35_2 & new_n3338_;
  assign new_n3340_ = ~new_n3335_ & ~new_n3339_;
  assign new_n3341_ = controlPi_35_4 & ~new_n3340_;
  assign new_n3342_ = controlPi_35_1 & n457_ntk1;
  assign new_n3343_ = ~controlPi_35_1 & n454_ntk1;
  assign new_n3344_ = ~new_n3342_ & ~new_n3343_;
  assign new_n3345_ = ~controlPi_35_2 & new_n3344_;
  assign new_n3346_ = controlPi_35_1 & n507_ntk1;
  assign new_n3347_ = ~controlPi_35_1 & n468_ntk1;
  assign new_n3348_ = ~new_n3346_ & ~new_n3347_;
  assign new_n3349_ = controlPi_35_2 & new_n3348_;
  assign new_n3350_ = ~new_n3345_ & ~new_n3349_;
  assign new_n3351_ = ~controlPi_35_4 & ~new_n3350_;
  assign new_n3352_ = ~new_n3341_ & ~new_n3351_;
  assign new_n3353_ = ~controlPi_35_3 & ~new_n3352_;
  assign new_n3354_ = controlPi_35_1 & n600_ntk1;
  assign new_n3355_ = ~controlPi_35_1 & n582_ntk1;
  assign new_n3356_ = ~new_n3354_ & ~new_n3355_;
  assign new_n3357_ = controlPi_35_2 & new_n3356_;
  assign new_n3358_ = controlPi_35_1 & n525_ntk1;
  assign new_n3359_ = ~controlPi_35_1 & n511_ntk1;
  assign new_n3360_ = ~new_n3358_ & ~new_n3359_;
  assign new_n3361_ = ~controlPi_35_2 & new_n3360_;
  assign new_n3362_ = ~new_n3357_ & ~new_n3361_;
  assign new_n3363_ = controlPi_35_3 & ~new_n3362_;
  assign new_n3364_ = ~controlPi_35_4 & new_n3363_;
  assign new_n3365_ = ~new_n3353_ & ~new_n3364_;
  assign new_n3366_ = controlPi_35_5 & ~new_n3365_;
  assign new_n3367_ = ~new_n3331_ & ~new_n3366_;
  assign new_n3368_ = controlPi_35_0 & ~new_n3367_;
  assign new_n3369_ = ~controlPi_35_0 & new_n3367_;
  assign new_n3370_ = ~new_n3368_ & ~new_n3369_;
  assign new_n3371_ = new_n2432_ & new_n3370_;
  assign new_n3372_ = new_n1946_ & new_n2689_;
  assign new_n3373_ = ~new_n2690_ & ~new_n3372_;
  assign new_n3374_ = ~new_n2432_ & ~new_n3373_;
  assign new_n3375_ = ~new_n3371_ & ~new_n3374_;
  assign new_n3376_ = new_n2146_ & ~new_n3375_;
  assign new_n3377_ = new_n1946_ & new_n2317_;
  assign new_n3378_ = ~new_n2318_ & ~new_n3377_;
  assign new_n3379_ = ~new_n2146_ & ~new_n3378_;
  assign new_n3380_ = ~new_n3376_ & ~new_n3379_;
  assign new_n3381_ = new_n1605_ & ~new_n3380_;
  assign new_n3382_ = ~new_n3285_ & ~new_n3381_;
  assign new_n3383_ = new_n1586_ & ~new_n3382_;
  assign new_n3384_ = ~new_n3282_ & ~new_n3383_;
  assign new_n3385_ = new_n1567_ & ~new_n3384_;
  assign new_n3386_ = new_n1281_ & ~new_n1567_;
  assign new_n3387_ = ~new_n3385_ & ~new_n3386_;
  assign new_n3388_ = ~new_n3281_ & new_n3387_;
  assign new_n3389_ = ~new_n3191_ & new_n3388_;
  assign new_n3390_ = new_n3075_ & ~new_n3389_;
  assign new_n3391_ = new_n3191_ & ~new_n3388_;
  assign new_n3392_ = ~new_n3390_ & ~new_n3391_;
  assign new_n3393_ = new_n939_ & ~new_n3392_;
  assign new_n3394_ = ~new_n3075_ & new_n3191_;
  assign new_n3395_ = new_n3075_ & ~new_n3191_;
  assign new_n3396_ = new_n3281_ & new_n3387_;
  assign new_n3397_ = ~new_n3395_ & ~new_n3396_;
  assign new_n3398_ = ~new_n3394_ & ~new_n3397_;
  assign new_n3399_ = ~new_n939_ & ~new_n3398_;
  assign new_n3400_ = ~new_n3393_ & ~new_n3399_;
  assign new_n3401_ = new_n2983_ & ~new_n3400_;
  assign new_n3402_ = ~new_n2983_ & new_n3400_;
  assign new_n3403_ = ~new_n3401_ & ~new_n3402_;
  assign new_n3404_ = new_n920_ & new_n3403_;
  assign new_n3405_ = ~new_n920_ & ~new_n3403_;
  assign new_n3406_ = ~n266_ntk1 & new_n870_;
  assign new_n3407_ = ~new_n865_ & ~new_n868_;
  assign new_n3408_ = ~new_n3406_ & new_n3407_;
  assign new_n3409_ = ~new_n911_ & ~new_n912_;
  assign new_n3410_ = new_n3408_ & new_n3409_;
  assign new_n3411_ = ~new_n3408_ & ~new_n3409_;
  assign new_n3412_ = ~new_n3410_ & ~new_n3411_;
  assign new_n3413_ = ~new_n3394_ & ~new_n3395_;
  assign new_n3414_ = new_n939_ & new_n3388_;
  assign new_n3415_ = ~new_n939_ & new_n3396_;
  assign new_n3416_ = ~new_n3414_ & ~new_n3415_;
  assign new_n3417_ = new_n3413_ & ~new_n3416_;
  assign new_n3418_ = ~new_n3413_ & new_n3416_;
  assign new_n3419_ = ~new_n3417_ & ~new_n3418_;
  assign new_n3420_ = new_n3412_ & new_n3419_;
  assign new_n3421_ = ~new_n3412_ & ~new_n3419_;
  assign new_n3422_ = new_n865_ & new_n870_;
  assign new_n3423_ = ~new_n913_ & ~new_n3422_;
  assign new_n3424_ = ~new_n3281_ & ~new_n3387_;
  assign new_n3425_ = ~new_n3396_ & ~new_n3424_;
  assign new_n3426_ = ~new_n3423_ & ~new_n3425_;
  assign new_n3427_ = new_n3423_ & new_n3425_;
  assign new_n3428_ = ~new_n3426_ & ~new_n3427_;
  assign new_n3429_ = ~new_n3421_ & new_n3428_;
  assign new_n3430_ = ~new_n3420_ & new_n3429_;
  assign new_n3431_ = ~new_n3405_ & new_n3430_;
  assign new_n3432_ = ~new_n3404_ & new_n3431_;
  assign new_n3433_ = n468_ntk1 & ~new_n825_;
  assign new_n3434_ = ~n468_ntk1 & new_n825_;
  assign new_n3435_ = ~new_n3433_ & ~new_n3434_;
  assign new_n3436_ = n616_ntk1 & new_n3435_;
  assign new_n3437_ = ~n616_ntk1 & ~new_n3435_;
  assign new_n3438_ = ~new_n3436_ & ~new_n3437_;
  assign new_n3439_ = ~new_n824_ & ~new_n828_;
  assign new_n3440_ = ~new_n829_ & ~new_n3439_;
  assign new_n3441_ = new_n3438_ & ~new_n3440_;
  assign new_n3442_ = ~new_n3438_ & new_n3440_;
  assign new_n3443_ = ~new_n3441_ & ~new_n3442_;
  assign new_n3444_ = n93_ntk1 & ~new_n3443_;
  assign new_n3445_ = new_n777_ & ~new_n779_;
  assign new_n3446_ = n349_ntk1 & ~new_n3445_;
  assign new_n3447_ = ~new_n778_ & new_n3446_;
  assign new_n3448_ = n199_ntk1 & new_n798_;
  assign new_n3449_ = new_n789_ & ~new_n791_;
  assign new_n3450_ = ~new_n790_ & new_n794_;
  assign new_n3451_ = ~new_n3449_ & new_n3450_;
  assign new_n3452_ = ~new_n3448_ & ~new_n3451_;
  assign new_n3453_ = ~new_n3447_ & new_n3452_;
  assign new_n3454_ = new_n772_ & ~new_n3453_;
  assign new_n3455_ = ~n616_ntk1 & ~new_n805_;
  assign new_n3456_ = n616_ntk1 & new_n805_;
  assign new_n3457_ = n206_ntk1 & ~new_n3456_;
  assign new_n3458_ = ~new_n3455_ & new_n3457_;
  assign new_n3459_ = new_n812_ & ~new_n814_;
  assign new_n3460_ = ~new_n813_ & new_n817_;
  assign new_n3461_ = ~new_n3459_ & new_n3460_;
  assign new_n3462_ = ~new_n3458_ & ~new_n3461_;
  assign new_n3463_ = ~new_n3454_ & new_n3462_;
  assign new_n3464_ = ~n93_ntk1 & ~new_n3463_;
  assign new_n3465_ = ~new_n3444_ & ~new_n3464_;
  assign new_n3466_ = ~n616_ntk1 & ~new_n839_;
  assign new_n3467_ = n616_ntk1 & new_n839_;
  assign new_n3468_ = ~new_n3466_ & ~new_n3467_;
  assign new_n3469_ = n266_ntk1 & ~new_n3468_;
  assign new_n3470_ = ~n266_ntk1 & ~n507_ntk1;
  assign new_n3471_ = ~new_n3469_ & ~new_n3470_;
  assign new_n3472_ = ~new_n3465_ & ~new_n3471_;
  assign new_n3473_ = new_n3465_ & new_n3471_;
  assign new_n3474_ = ~new_n3472_ & ~new_n3473_;
  assign new_n3475_ = ~new_n844_ & ~new_n909_;
  assign new_n3476_ = ~new_n845_ & ~new_n3475_;
  assign new_n3477_ = n266_ntk1 & new_n3476_;
  assign new_n3478_ = ~new_n843_ & new_n915_;
  assign new_n3479_ = ~new_n835_ & ~new_n3478_;
  assign new_n3480_ = new_n843_ & ~new_n915_;
  assign new_n3481_ = ~new_n3479_ & ~new_n3480_;
  assign new_n3482_ = ~n266_ntk1 & ~new_n3481_;
  assign new_n3483_ = ~new_n3477_ & ~new_n3482_;
  assign new_n3484_ = new_n3474_ & new_n3483_;
  assign new_n3485_ = ~new_n3474_ & ~new_n3483_;
  assign new_n3486_ = ~new_n3484_ & ~new_n3485_;
  assign new_n3487_ = ~controlPi_34_1 & ~n199_ntk1;
  assign new_n3488_ = controlPi_34_1 & ~n211_ntk1;
  assign new_n3489_ = ~new_n3487_ & ~new_n3488_;
  assign new_n3490_ = ~controlPi_34_2 & new_n3489_;
  assign new_n3491_ = ~controlPi_34_1 & ~n216_ntk1;
  assign new_n3492_ = controlPi_34_1 & ~n280_ntk1;
  assign new_n3493_ = ~new_n3491_ & ~new_n3492_;
  assign new_n3494_ = controlPi_34_2 & new_n3493_;
  assign new_n3495_ = ~new_n3490_ & ~new_n3494_;
  assign new_n3496_ = ~controlPi_34_3 & new_n3495_;
  assign new_n3497_ = ~controlPi_34_1 & ~n287_ntk1;
  assign new_n3498_ = controlPi_34_1 & ~n409_ntk1;
  assign new_n3499_ = ~new_n3497_ & ~new_n3498_;
  assign new_n3500_ = ~controlPi_34_2 & new_n3499_;
  assign new_n3501_ = ~controlPi_34_1 & ~n428_ntk1;
  assign new_n3502_ = controlPi_34_1 & ~n435_ntk1;
  assign new_n3503_ = ~new_n3501_ & ~new_n3502_;
  assign new_n3504_ = controlPi_34_2 & new_n3503_;
  assign new_n3505_ = ~new_n3500_ & ~new_n3504_;
  assign new_n3506_ = controlPi_34_3 & new_n3505_;
  assign new_n3507_ = ~new_n3496_ & ~new_n3506_;
  assign new_n3508_ = controlPi_34_4 & ~new_n3507_;
  assign new_n3509_ = ~controlPi_34_1 & ~n2_ntk1;
  assign new_n3510_ = controlPi_34_1 & ~n13_ntk1;
  assign new_n3511_ = ~new_n3509_ & ~new_n3510_;
  assign new_n3512_ = ~controlPi_34_2 & new_n3511_;
  assign new_n3513_ = ~controlPi_34_1 & ~n46_ntk1;
  assign new_n3514_ = controlPi_34_1 & ~n75_ntk1;
  assign new_n3515_ = ~new_n3513_ & ~new_n3514_;
  assign new_n3516_ = controlPi_34_2 & new_n3515_;
  assign new_n3517_ = ~new_n3512_ & ~new_n3516_;
  assign new_n3518_ = ~controlPi_34_3 & new_n3517_;
  assign new_n3519_ = ~controlPi_34_1 & ~n96_ntk1;
  assign new_n3520_ = controlPi_34_1 & ~n131_ntk1;
  assign new_n3521_ = ~new_n3519_ & ~new_n3520_;
  assign new_n3522_ = ~controlPi_34_2 & new_n3521_;
  assign new_n3523_ = ~controlPi_34_1 & ~n159_ntk1;
  assign new_n3524_ = controlPi_34_1 & ~n177_ntk1;
  assign new_n3525_ = ~new_n3523_ & ~new_n3524_;
  assign new_n3526_ = controlPi_34_2 & new_n3525_;
  assign new_n3527_ = ~new_n3522_ & ~new_n3526_;
  assign new_n3528_ = controlPi_34_3 & new_n3527_;
  assign new_n3529_ = ~new_n3518_ & ~new_n3528_;
  assign new_n3530_ = ~controlPi_34_4 & ~new_n3529_;
  assign new_n3531_ = ~new_n3508_ & ~new_n3530_;
  assign new_n3532_ = ~controlPi_34_5 & ~new_n3531_;
  assign new_n3533_ = controlPi_34_1 & n659_ntk1;
  assign new_n3534_ = ~controlPi_34_1 & n616_ntk1;
  assign new_n3535_ = ~new_n3533_ & ~new_n3534_;
  assign new_n3536_ = ~controlPi_34_2 & new_n3535_;
  assign new_n3537_ = controlPi_34_1 & n673_ntk1;
  assign new_n3538_ = ~controlPi_34_1 & n664_ntk1;
  assign new_n3539_ = ~new_n3537_ & ~new_n3538_;
  assign new_n3540_ = controlPi_34_2 & new_n3539_;
  assign new_n3541_ = ~new_n3536_ & ~new_n3540_;
  assign new_n3542_ = controlPi_34_4 & ~new_n3541_;
  assign new_n3543_ = controlPi_34_1 & n457_ntk1;
  assign new_n3544_ = ~controlPi_34_1 & n454_ntk1;
  assign new_n3545_ = ~new_n3543_ & ~new_n3544_;
  assign new_n3546_ = ~controlPi_34_2 & new_n3545_;
  assign new_n3547_ = controlPi_34_1 & n507_ntk1;
  assign new_n3548_ = ~controlPi_34_1 & n468_ntk1;
  assign new_n3549_ = ~new_n3547_ & ~new_n3548_;
  assign new_n3550_ = controlPi_34_2 & new_n3549_;
  assign new_n3551_ = ~new_n3546_ & ~new_n3550_;
  assign new_n3552_ = ~controlPi_34_4 & ~new_n3551_;
  assign new_n3553_ = ~new_n3542_ & ~new_n3552_;
  assign new_n3554_ = ~controlPi_34_3 & ~new_n3553_;
  assign new_n3555_ = controlPi_34_1 & n600_ntk1;
  assign new_n3556_ = ~controlPi_34_1 & n582_ntk1;
  assign new_n3557_ = ~new_n3555_ & ~new_n3556_;
  assign new_n3558_ = controlPi_34_2 & new_n3557_;
  assign new_n3559_ = controlPi_34_1 & n525_ntk1;
  assign new_n3560_ = ~controlPi_34_1 & n511_ntk1;
  assign new_n3561_ = ~new_n3559_ & ~new_n3560_;
  assign new_n3562_ = ~controlPi_34_2 & new_n3561_;
  assign new_n3563_ = ~new_n3558_ & ~new_n3562_;
  assign new_n3564_ = controlPi_34_3 & ~new_n3563_;
  assign new_n3565_ = ~controlPi_34_4 & new_n3564_;
  assign new_n3566_ = ~new_n3554_ & ~new_n3565_;
  assign new_n3567_ = controlPi_34_5 & ~new_n3566_;
  assign new_n3568_ = ~new_n3532_ & ~new_n3567_;
  assign new_n3569_ = controlPi_34_0 & ~new_n3568_;
  assign new_n3570_ = ~controlPi_34_0 & new_n3568_;
  assign new_n3571_ = ~new_n3569_ & ~new_n3570_;
  assign new_n3572_ = new_n939_ & ~new_n3571_;
  assign new_n3573_ = ~new_n1370_ & ~new_n1542_;
  assign new_n3574_ = ~new_n1541_ & ~new_n3573_;
  assign new_n3575_ = ~controlPi_19_1 & ~n199_ntk1;
  assign new_n3576_ = controlPi_19_1 & ~n211_ntk1;
  assign new_n3577_ = ~new_n3575_ & ~new_n3576_;
  assign new_n3578_ = ~controlPi_19_2 & new_n3577_;
  assign new_n3579_ = ~controlPi_19_1 & ~n216_ntk1;
  assign new_n3580_ = controlPi_19_1 & ~n280_ntk1;
  assign new_n3581_ = ~new_n3579_ & ~new_n3580_;
  assign new_n3582_ = controlPi_19_2 & new_n3581_;
  assign new_n3583_ = ~new_n3578_ & ~new_n3582_;
  assign new_n3584_ = ~controlPi_19_3 & new_n3583_;
  assign new_n3585_ = ~controlPi_19_1 & ~n287_ntk1;
  assign new_n3586_ = controlPi_19_1 & ~n409_ntk1;
  assign new_n3587_ = ~new_n3585_ & ~new_n3586_;
  assign new_n3588_ = ~controlPi_19_2 & new_n3587_;
  assign new_n3589_ = ~controlPi_19_1 & ~n428_ntk1;
  assign new_n3590_ = controlPi_19_1 & ~n435_ntk1;
  assign new_n3591_ = ~new_n3589_ & ~new_n3590_;
  assign new_n3592_ = controlPi_19_2 & new_n3591_;
  assign new_n3593_ = ~new_n3588_ & ~new_n3592_;
  assign new_n3594_ = controlPi_19_3 & new_n3593_;
  assign new_n3595_ = ~new_n3584_ & ~new_n3594_;
  assign new_n3596_ = controlPi_19_4 & ~new_n3595_;
  assign new_n3597_ = ~controlPi_19_1 & ~n2_ntk1;
  assign new_n3598_ = controlPi_19_1 & ~n13_ntk1;
  assign new_n3599_ = ~new_n3597_ & ~new_n3598_;
  assign new_n3600_ = ~controlPi_19_2 & new_n3599_;
  assign new_n3601_ = ~controlPi_19_1 & ~n46_ntk1;
  assign new_n3602_ = controlPi_19_1 & ~n75_ntk1;
  assign new_n3603_ = ~new_n3601_ & ~new_n3602_;
  assign new_n3604_ = controlPi_19_2 & new_n3603_;
  assign new_n3605_ = ~new_n3600_ & ~new_n3604_;
  assign new_n3606_ = ~controlPi_19_3 & new_n3605_;
  assign new_n3607_ = ~controlPi_19_1 & ~n96_ntk1;
  assign new_n3608_ = controlPi_19_1 & ~n131_ntk1;
  assign new_n3609_ = ~new_n3607_ & ~new_n3608_;
  assign new_n3610_ = ~controlPi_19_2 & new_n3609_;
  assign new_n3611_ = ~controlPi_19_1 & ~n159_ntk1;
  assign new_n3612_ = controlPi_19_1 & ~n177_ntk1;
  assign new_n3613_ = ~new_n3611_ & ~new_n3612_;
  assign new_n3614_ = controlPi_19_2 & new_n3613_;
  assign new_n3615_ = ~new_n3610_ & ~new_n3614_;
  assign new_n3616_ = controlPi_19_3 & new_n3615_;
  assign new_n3617_ = ~new_n3606_ & ~new_n3616_;
  assign new_n3618_ = ~controlPi_19_4 & ~new_n3617_;
  assign new_n3619_ = ~new_n3596_ & ~new_n3618_;
  assign new_n3620_ = ~controlPi_19_5 & ~new_n3619_;
  assign new_n3621_ = controlPi_19_1 & n659_ntk1;
  assign new_n3622_ = ~controlPi_19_1 & n616_ntk1;
  assign new_n3623_ = ~new_n3621_ & ~new_n3622_;
  assign new_n3624_ = ~controlPi_19_2 & new_n3623_;
  assign new_n3625_ = controlPi_19_1 & n673_ntk1;
  assign new_n3626_ = ~controlPi_19_1 & n664_ntk1;
  assign new_n3627_ = ~new_n3625_ & ~new_n3626_;
  assign new_n3628_ = controlPi_19_2 & new_n3627_;
  assign new_n3629_ = ~new_n3624_ & ~new_n3628_;
  assign new_n3630_ = controlPi_19_4 & ~new_n3629_;
  assign new_n3631_ = controlPi_19_1 & n457_ntk1;
  assign new_n3632_ = ~controlPi_19_1 & n454_ntk1;
  assign new_n3633_ = ~new_n3631_ & ~new_n3632_;
  assign new_n3634_ = ~controlPi_19_2 & new_n3633_;
  assign new_n3635_ = controlPi_19_1 & n507_ntk1;
  assign new_n3636_ = ~controlPi_19_1 & n468_ntk1;
  assign new_n3637_ = ~new_n3635_ & ~new_n3636_;
  assign new_n3638_ = controlPi_19_2 & new_n3637_;
  assign new_n3639_ = ~new_n3634_ & ~new_n3638_;
  assign new_n3640_ = ~controlPi_19_4 & ~new_n3639_;
  assign new_n3641_ = ~new_n3630_ & ~new_n3640_;
  assign new_n3642_ = ~controlPi_19_3 & ~new_n3641_;
  assign new_n3643_ = controlPi_19_1 & n600_ntk1;
  assign new_n3644_ = ~controlPi_19_1 & n582_ntk1;
  assign new_n3645_ = ~new_n3643_ & ~new_n3644_;
  assign new_n3646_ = controlPi_19_2 & new_n3645_;
  assign new_n3647_ = controlPi_19_1 & n525_ntk1;
  assign new_n3648_ = ~controlPi_19_1 & n511_ntk1;
  assign new_n3649_ = ~new_n3647_ & ~new_n3648_;
  assign new_n3650_ = ~controlPi_19_2 & new_n3649_;
  assign new_n3651_ = ~new_n3646_ & ~new_n3650_;
  assign new_n3652_ = controlPi_19_3 & ~new_n3651_;
  assign new_n3653_ = ~controlPi_19_4 & new_n3652_;
  assign new_n3654_ = ~new_n3642_ & ~new_n3653_;
  assign new_n3655_ = controlPi_19_5 & ~new_n3654_;
  assign new_n3656_ = ~new_n3620_ & ~new_n3655_;
  assign new_n3657_ = controlPi_19_0 & ~new_n3656_;
  assign new_n3658_ = ~controlPi_19_0 & new_n3656_;
  assign new_n3659_ = ~new_n3657_ & ~new_n3658_;
  assign new_n3660_ = ~controlPi_54_1 & ~n199_ntk1;
  assign new_n3661_ = controlPi_54_1 & ~n211_ntk1;
  assign new_n3662_ = ~new_n3660_ & ~new_n3661_;
  assign new_n3663_ = ~controlPi_54_2 & new_n3662_;
  assign new_n3664_ = ~controlPi_54_1 & ~n216_ntk1;
  assign new_n3665_ = controlPi_54_1 & ~n280_ntk1;
  assign new_n3666_ = ~new_n3664_ & ~new_n3665_;
  assign new_n3667_ = controlPi_54_2 & new_n3666_;
  assign new_n3668_ = ~new_n3663_ & ~new_n3667_;
  assign new_n3669_ = ~controlPi_54_3 & new_n3668_;
  assign new_n3670_ = ~controlPi_54_1 & ~n287_ntk1;
  assign new_n3671_ = controlPi_54_1 & ~n409_ntk1;
  assign new_n3672_ = ~new_n3670_ & ~new_n3671_;
  assign new_n3673_ = ~controlPi_54_2 & new_n3672_;
  assign new_n3674_ = ~controlPi_54_1 & ~n428_ntk1;
  assign new_n3675_ = controlPi_54_1 & ~n435_ntk1;
  assign new_n3676_ = ~new_n3674_ & ~new_n3675_;
  assign new_n3677_ = controlPi_54_2 & new_n3676_;
  assign new_n3678_ = ~new_n3673_ & ~new_n3677_;
  assign new_n3679_ = controlPi_54_3 & new_n3678_;
  assign new_n3680_ = ~new_n3669_ & ~new_n3679_;
  assign new_n3681_ = controlPi_54_4 & ~new_n3680_;
  assign new_n3682_ = ~controlPi_54_1 & ~n2_ntk1;
  assign new_n3683_ = controlPi_54_1 & ~n13_ntk1;
  assign new_n3684_ = ~new_n3682_ & ~new_n3683_;
  assign new_n3685_ = ~controlPi_54_2 & new_n3684_;
  assign new_n3686_ = ~controlPi_54_1 & ~n46_ntk1;
  assign new_n3687_ = controlPi_54_1 & ~n75_ntk1;
  assign new_n3688_ = ~new_n3686_ & ~new_n3687_;
  assign new_n3689_ = controlPi_54_2 & new_n3688_;
  assign new_n3690_ = ~new_n3685_ & ~new_n3689_;
  assign new_n3691_ = ~controlPi_54_3 & new_n3690_;
  assign new_n3692_ = ~controlPi_54_1 & ~n96_ntk1;
  assign new_n3693_ = controlPi_54_1 & ~n131_ntk1;
  assign new_n3694_ = ~new_n3692_ & ~new_n3693_;
  assign new_n3695_ = ~controlPi_54_2 & new_n3694_;
  assign new_n3696_ = ~controlPi_54_1 & ~n159_ntk1;
  assign new_n3697_ = controlPi_54_1 & ~n177_ntk1;
  assign new_n3698_ = ~new_n3696_ & ~new_n3697_;
  assign new_n3699_ = controlPi_54_2 & new_n3698_;
  assign new_n3700_ = ~new_n3695_ & ~new_n3699_;
  assign new_n3701_ = controlPi_54_3 & new_n3700_;
  assign new_n3702_ = ~new_n3691_ & ~new_n3701_;
  assign new_n3703_ = ~controlPi_54_4 & ~new_n3702_;
  assign new_n3704_ = ~new_n3681_ & ~new_n3703_;
  assign new_n3705_ = ~controlPi_54_5 & ~new_n3704_;
  assign new_n3706_ = controlPi_54_1 & n659_ntk1;
  assign new_n3707_ = ~controlPi_54_1 & n616_ntk1;
  assign new_n3708_ = ~new_n3706_ & ~new_n3707_;
  assign new_n3709_ = ~controlPi_54_2 & new_n3708_;
  assign new_n3710_ = controlPi_54_1 & n673_ntk1;
  assign new_n3711_ = ~controlPi_54_1 & n664_ntk1;
  assign new_n3712_ = ~new_n3710_ & ~new_n3711_;
  assign new_n3713_ = controlPi_54_2 & new_n3712_;
  assign new_n3714_ = ~new_n3709_ & ~new_n3713_;
  assign new_n3715_ = controlPi_54_4 & ~new_n3714_;
  assign new_n3716_ = controlPi_54_1 & n457_ntk1;
  assign new_n3717_ = ~controlPi_54_1 & n454_ntk1;
  assign new_n3718_ = ~new_n3716_ & ~new_n3717_;
  assign new_n3719_ = ~controlPi_54_2 & new_n3718_;
  assign new_n3720_ = controlPi_54_1 & n507_ntk1;
  assign new_n3721_ = ~controlPi_54_1 & n468_ntk1;
  assign new_n3722_ = ~new_n3720_ & ~new_n3721_;
  assign new_n3723_ = controlPi_54_2 & new_n3722_;
  assign new_n3724_ = ~new_n3719_ & ~new_n3723_;
  assign new_n3725_ = ~controlPi_54_4 & ~new_n3724_;
  assign new_n3726_ = ~new_n3715_ & ~new_n3725_;
  assign new_n3727_ = ~controlPi_54_3 & ~new_n3726_;
  assign new_n3728_ = controlPi_54_1 & n600_ntk1;
  assign new_n3729_ = ~controlPi_54_1 & n582_ntk1;
  assign new_n3730_ = ~new_n3728_ & ~new_n3729_;
  assign new_n3731_ = controlPi_54_2 & new_n3730_;
  assign new_n3732_ = controlPi_54_1 & n525_ntk1;
  assign new_n3733_ = ~controlPi_54_1 & n511_ntk1;
  assign new_n3734_ = ~new_n3732_ & ~new_n3733_;
  assign new_n3735_ = ~controlPi_54_2 & new_n3734_;
  assign new_n3736_ = ~new_n3731_ & ~new_n3735_;
  assign new_n3737_ = controlPi_54_3 & ~new_n3736_;
  assign new_n3738_ = ~controlPi_54_4 & new_n3737_;
  assign new_n3739_ = ~new_n3727_ & ~new_n3738_;
  assign new_n3740_ = controlPi_54_5 & ~new_n3739_;
  assign new_n3741_ = ~new_n3705_ & ~new_n3740_;
  assign new_n3742_ = controlPi_54_0 & ~new_n3741_;
  assign new_n3743_ = ~controlPi_54_0 & new_n3741_;
  assign new_n3744_ = ~new_n3742_ & ~new_n3743_;
  assign new_n3745_ = ~new_n3659_ & new_n3744_;
  assign new_n3746_ = new_n3659_ & ~new_n3744_;
  assign new_n3747_ = ~new_n3745_ & ~new_n3746_;
  assign new_n3748_ = new_n3574_ & new_n3747_;
  assign new_n3749_ = ~new_n3574_ & ~new_n3747_;
  assign new_n3750_ = ~new_n939_ & ~new_n3749_;
  assign new_n3751_ = ~new_n3748_ & new_n3750_;
  assign new_n3752_ = ~new_n3572_ & ~new_n3751_;
  assign new_n3753_ = ~new_n2971_ & ~new_n2974_;
  assign new_n3754_ = ~new_n2973_ & ~new_n3753_;
  assign new_n3755_ = ~controlPi_73_1 & ~n199_ntk1;
  assign new_n3756_ = controlPi_73_1 & ~n211_ntk1;
  assign new_n3757_ = ~new_n3755_ & ~new_n3756_;
  assign new_n3758_ = ~controlPi_73_2 & new_n3757_;
  assign new_n3759_ = ~controlPi_73_1 & ~n216_ntk1;
  assign new_n3760_ = controlPi_73_1 & ~n280_ntk1;
  assign new_n3761_ = ~new_n3759_ & ~new_n3760_;
  assign new_n3762_ = controlPi_73_2 & new_n3761_;
  assign new_n3763_ = ~new_n3758_ & ~new_n3762_;
  assign new_n3764_ = ~controlPi_73_3 & new_n3763_;
  assign new_n3765_ = ~controlPi_73_1 & ~n287_ntk1;
  assign new_n3766_ = controlPi_73_1 & ~n409_ntk1;
  assign new_n3767_ = ~new_n3765_ & ~new_n3766_;
  assign new_n3768_ = ~controlPi_73_2 & new_n3767_;
  assign new_n3769_ = ~controlPi_73_1 & ~n428_ntk1;
  assign new_n3770_ = controlPi_73_1 & ~n435_ntk1;
  assign new_n3771_ = ~new_n3769_ & ~new_n3770_;
  assign new_n3772_ = controlPi_73_2 & new_n3771_;
  assign new_n3773_ = ~new_n3768_ & ~new_n3772_;
  assign new_n3774_ = controlPi_73_3 & new_n3773_;
  assign new_n3775_ = ~new_n3764_ & ~new_n3774_;
  assign new_n3776_ = controlPi_73_4 & ~new_n3775_;
  assign new_n3777_ = ~controlPi_73_1 & ~n2_ntk1;
  assign new_n3778_ = controlPi_73_1 & ~n13_ntk1;
  assign new_n3779_ = ~new_n3777_ & ~new_n3778_;
  assign new_n3780_ = ~controlPi_73_2 & new_n3779_;
  assign new_n3781_ = ~controlPi_73_1 & ~n46_ntk1;
  assign new_n3782_ = controlPi_73_1 & ~n75_ntk1;
  assign new_n3783_ = ~new_n3781_ & ~new_n3782_;
  assign new_n3784_ = controlPi_73_2 & new_n3783_;
  assign new_n3785_ = ~new_n3780_ & ~new_n3784_;
  assign new_n3786_ = ~controlPi_73_3 & new_n3785_;
  assign new_n3787_ = ~controlPi_73_1 & ~n96_ntk1;
  assign new_n3788_ = controlPi_73_1 & ~n131_ntk1;
  assign new_n3789_ = ~new_n3787_ & ~new_n3788_;
  assign new_n3790_ = ~controlPi_73_2 & new_n3789_;
  assign new_n3791_ = ~controlPi_73_1 & ~n159_ntk1;
  assign new_n3792_ = controlPi_73_1 & ~n177_ntk1;
  assign new_n3793_ = ~new_n3791_ & ~new_n3792_;
  assign new_n3794_ = controlPi_73_2 & new_n3793_;
  assign new_n3795_ = ~new_n3790_ & ~new_n3794_;
  assign new_n3796_ = controlPi_73_3 & new_n3795_;
  assign new_n3797_ = ~new_n3786_ & ~new_n3796_;
  assign new_n3798_ = ~controlPi_73_4 & ~new_n3797_;
  assign new_n3799_ = ~new_n3776_ & ~new_n3798_;
  assign new_n3800_ = ~controlPi_73_5 & ~new_n3799_;
  assign new_n3801_ = controlPi_73_1 & n659_ntk1;
  assign new_n3802_ = ~controlPi_73_1 & n616_ntk1;
  assign new_n3803_ = ~new_n3801_ & ~new_n3802_;
  assign new_n3804_ = ~controlPi_73_2 & new_n3803_;
  assign new_n3805_ = controlPi_73_1 & n673_ntk1;
  assign new_n3806_ = ~controlPi_73_1 & n664_ntk1;
  assign new_n3807_ = ~new_n3805_ & ~new_n3806_;
  assign new_n3808_ = controlPi_73_2 & new_n3807_;
  assign new_n3809_ = ~new_n3804_ & ~new_n3808_;
  assign new_n3810_ = controlPi_73_4 & ~new_n3809_;
  assign new_n3811_ = controlPi_73_1 & n457_ntk1;
  assign new_n3812_ = ~controlPi_73_1 & n454_ntk1;
  assign new_n3813_ = ~new_n3811_ & ~new_n3812_;
  assign new_n3814_ = ~controlPi_73_2 & new_n3813_;
  assign new_n3815_ = controlPi_73_1 & n507_ntk1;
  assign new_n3816_ = ~controlPi_73_1 & n468_ntk1;
  assign new_n3817_ = ~new_n3815_ & ~new_n3816_;
  assign new_n3818_ = controlPi_73_2 & new_n3817_;
  assign new_n3819_ = ~new_n3814_ & ~new_n3818_;
  assign new_n3820_ = ~controlPi_73_4 & ~new_n3819_;
  assign new_n3821_ = ~new_n3810_ & ~new_n3820_;
  assign new_n3822_ = ~controlPi_73_3 & ~new_n3821_;
  assign new_n3823_ = controlPi_73_1 & n600_ntk1;
  assign new_n3824_ = ~controlPi_73_1 & n582_ntk1;
  assign new_n3825_ = ~new_n3823_ & ~new_n3824_;
  assign new_n3826_ = controlPi_73_2 & new_n3825_;
  assign new_n3827_ = controlPi_73_1 & n525_ntk1;
  assign new_n3828_ = ~controlPi_73_1 & n511_ntk1;
  assign new_n3829_ = ~new_n3827_ & ~new_n3828_;
  assign new_n3830_ = ~controlPi_73_2 & new_n3829_;
  assign new_n3831_ = ~new_n3826_ & ~new_n3830_;
  assign new_n3832_ = controlPi_73_3 & ~new_n3831_;
  assign new_n3833_ = ~controlPi_73_4 & new_n3832_;
  assign new_n3834_ = ~new_n3822_ & ~new_n3833_;
  assign new_n3835_ = controlPi_73_5 & ~new_n3834_;
  assign new_n3836_ = ~new_n3800_ & ~new_n3835_;
  assign new_n3837_ = controlPi_73_0 & ~new_n3836_;
  assign new_n3838_ = ~controlPi_73_0 & new_n3836_;
  assign new_n3839_ = ~new_n3837_ & ~new_n3838_;
  assign new_n3840_ = ~new_n2970_ & ~new_n3839_;
  assign new_n3841_ = new_n2970_ & new_n3839_;
  assign new_n3842_ = ~new_n3840_ & ~new_n3841_;
  assign new_n3843_ = ~new_n3744_ & ~new_n3842_;
  assign new_n3844_ = new_n3744_ & new_n3842_;
  assign new_n3845_ = ~new_n3843_ & ~new_n3844_;
  assign new_n3846_ = ~new_n3754_ & ~new_n3845_;
  assign new_n3847_ = new_n3754_ & new_n3845_;
  assign new_n3848_ = ~new_n3846_ & ~new_n3847_;
  assign new_n3849_ = ~new_n1567_ & ~new_n3848_;
  assign new_n3850_ = new_n1950_ & ~new_n2122_;
  assign new_n3851_ = ~new_n2121_ & ~new_n3850_;
  assign new_n3852_ = ~new_n1605_ & ~new_n3851_;
  assign new_n3853_ = new_n2321_ & ~new_n2408_;
  assign new_n3854_ = ~new_n2407_ & ~new_n3853_;
  assign new_n3855_ = ~new_n2146_ & ~new_n3854_;
  assign new_n3856_ = new_n2693_ & ~new_n2780_;
  assign new_n3857_ = ~new_n2779_ & ~new_n3856_;
  assign new_n3858_ = ~new_n2432_ & ~new_n3857_;
  assign new_n3859_ = ~controlPi_82_1 & ~n199_ntk1;
  assign new_n3860_ = controlPi_82_1 & ~n211_ntk1;
  assign new_n3861_ = ~new_n3859_ & ~new_n3860_;
  assign new_n3862_ = ~controlPi_82_2 & new_n3861_;
  assign new_n3863_ = ~controlPi_82_1 & ~n216_ntk1;
  assign new_n3864_ = controlPi_82_1 & ~n280_ntk1;
  assign new_n3865_ = ~new_n3863_ & ~new_n3864_;
  assign new_n3866_ = controlPi_82_2 & new_n3865_;
  assign new_n3867_ = ~new_n3862_ & ~new_n3866_;
  assign new_n3868_ = ~controlPi_82_3 & new_n3867_;
  assign new_n3869_ = ~controlPi_82_1 & ~n287_ntk1;
  assign new_n3870_ = controlPi_82_1 & ~n409_ntk1;
  assign new_n3871_ = ~new_n3869_ & ~new_n3870_;
  assign new_n3872_ = ~controlPi_82_2 & new_n3871_;
  assign new_n3873_ = ~controlPi_82_1 & ~n428_ntk1;
  assign new_n3874_ = controlPi_82_1 & ~n435_ntk1;
  assign new_n3875_ = ~new_n3873_ & ~new_n3874_;
  assign new_n3876_ = controlPi_82_2 & new_n3875_;
  assign new_n3877_ = ~new_n3872_ & ~new_n3876_;
  assign new_n3878_ = controlPi_82_3 & new_n3877_;
  assign new_n3879_ = ~new_n3868_ & ~new_n3878_;
  assign new_n3880_ = controlPi_82_4 & ~new_n3879_;
  assign new_n3881_ = ~controlPi_82_1 & ~n2_ntk1;
  assign new_n3882_ = controlPi_82_1 & ~n13_ntk1;
  assign new_n3883_ = ~new_n3881_ & ~new_n3882_;
  assign new_n3884_ = ~controlPi_82_2 & new_n3883_;
  assign new_n3885_ = ~controlPi_82_1 & ~n46_ntk1;
  assign new_n3886_ = controlPi_82_1 & ~n75_ntk1;
  assign new_n3887_ = ~new_n3885_ & ~new_n3886_;
  assign new_n3888_ = controlPi_82_2 & new_n3887_;
  assign new_n3889_ = ~new_n3884_ & ~new_n3888_;
  assign new_n3890_ = ~controlPi_82_3 & new_n3889_;
  assign new_n3891_ = ~controlPi_82_1 & ~n96_ntk1;
  assign new_n3892_ = controlPi_82_1 & ~n131_ntk1;
  assign new_n3893_ = ~new_n3891_ & ~new_n3892_;
  assign new_n3894_ = ~controlPi_82_2 & new_n3893_;
  assign new_n3895_ = ~controlPi_82_1 & ~n159_ntk1;
  assign new_n3896_ = controlPi_82_1 & ~n177_ntk1;
  assign new_n3897_ = ~new_n3895_ & ~new_n3896_;
  assign new_n3898_ = controlPi_82_2 & new_n3897_;
  assign new_n3899_ = ~new_n3894_ & ~new_n3898_;
  assign new_n3900_ = controlPi_82_3 & new_n3899_;
  assign new_n3901_ = ~new_n3890_ & ~new_n3900_;
  assign new_n3902_ = ~controlPi_82_4 & ~new_n3901_;
  assign new_n3903_ = ~new_n3880_ & ~new_n3902_;
  assign new_n3904_ = ~controlPi_82_5 & ~new_n3903_;
  assign new_n3905_ = controlPi_82_1 & n659_ntk1;
  assign new_n3906_ = ~controlPi_82_1 & n616_ntk1;
  assign new_n3907_ = ~new_n3905_ & ~new_n3906_;
  assign new_n3908_ = ~controlPi_82_2 & new_n3907_;
  assign new_n3909_ = controlPi_82_1 & n673_ntk1;
  assign new_n3910_ = ~controlPi_82_1 & n664_ntk1;
  assign new_n3911_ = ~new_n3909_ & ~new_n3910_;
  assign new_n3912_ = controlPi_82_2 & new_n3911_;
  assign new_n3913_ = ~new_n3908_ & ~new_n3912_;
  assign new_n3914_ = controlPi_82_4 & ~new_n3913_;
  assign new_n3915_ = controlPi_82_1 & n457_ntk1;
  assign new_n3916_ = ~controlPi_82_1 & n454_ntk1;
  assign new_n3917_ = ~new_n3915_ & ~new_n3916_;
  assign new_n3918_ = ~controlPi_82_2 & new_n3917_;
  assign new_n3919_ = controlPi_82_1 & n507_ntk1;
  assign new_n3920_ = ~controlPi_82_1 & n468_ntk1;
  assign new_n3921_ = ~new_n3919_ & ~new_n3920_;
  assign new_n3922_ = controlPi_82_2 & new_n3921_;
  assign new_n3923_ = ~new_n3918_ & ~new_n3922_;
  assign new_n3924_ = ~controlPi_82_4 & ~new_n3923_;
  assign new_n3925_ = ~new_n3914_ & ~new_n3924_;
  assign new_n3926_ = ~controlPi_82_3 & ~new_n3925_;
  assign new_n3927_ = controlPi_82_1 & n600_ntk1;
  assign new_n3928_ = ~controlPi_82_1 & n582_ntk1;
  assign new_n3929_ = ~new_n3927_ & ~new_n3928_;
  assign new_n3930_ = controlPi_82_2 & new_n3929_;
  assign new_n3931_ = controlPi_82_1 & n525_ntk1;
  assign new_n3932_ = ~controlPi_82_1 & n511_ntk1;
  assign new_n3933_ = ~new_n3931_ & ~new_n3932_;
  assign new_n3934_ = ~controlPi_82_2 & new_n3933_;
  assign new_n3935_ = ~new_n3930_ & ~new_n3934_;
  assign new_n3936_ = controlPi_82_3 & ~new_n3935_;
  assign new_n3937_ = ~controlPi_82_4 & new_n3936_;
  assign new_n3938_ = ~new_n3926_ & ~new_n3937_;
  assign new_n3939_ = controlPi_82_5 & ~new_n3938_;
  assign new_n3940_ = ~new_n3904_ & ~new_n3939_;
  assign new_n3941_ = ~controlPi_82_0 & ~new_n3940_;
  assign new_n3942_ = controlPi_82_0 & new_n3940_;
  assign new_n3943_ = ~new_n3941_ & ~new_n3942_;
  assign new_n3944_ = new_n2432_ & ~new_n3943_;
  assign new_n3945_ = ~new_n3858_ & ~new_n3944_;
  assign new_n3946_ = new_n2146_ & ~new_n3945_;
  assign new_n3947_ = ~new_n3855_ & ~new_n3946_;
  assign new_n3948_ = new_n1605_ & ~new_n3947_;
  assign new_n3949_ = ~new_n3852_ & ~new_n3948_;
  assign new_n3950_ = new_n1586_ & ~new_n3949_;
  assign new_n3951_ = ~new_n2794_ & ~new_n3744_;
  assign new_n3952_ = new_n2794_ & new_n3744_;
  assign new_n3953_ = ~new_n3951_ & ~new_n3952_;
  assign new_n3954_ = ~new_n1586_ & new_n3953_;
  assign new_n3955_ = ~new_n3950_ & ~new_n3954_;
  assign new_n3956_ = new_n1567_ & ~new_n3955_;
  assign new_n3957_ = ~new_n3849_ & ~new_n3956_;
  assign new_n3958_ = ~new_n3752_ & new_n3957_;
  assign new_n3959_ = new_n3752_ & ~new_n3957_;
  assign new_n3960_ = ~new_n3958_ & ~new_n3959_;
  assign new_n3961_ = ~new_n2982_ & ~new_n3398_;
  assign new_n3962_ = ~new_n2981_ & ~new_n3961_;
  assign new_n3963_ = ~new_n939_ & ~new_n3962_;
  assign new_n3964_ = new_n2980_ & new_n3392_;
  assign new_n3965_ = new_n1548_ & ~new_n3964_;
  assign new_n3966_ = ~new_n2980_ & ~new_n3392_;
  assign new_n3967_ = ~new_n3965_ & ~new_n3966_;
  assign new_n3968_ = new_n939_ & ~new_n3967_;
  assign new_n3969_ = ~new_n3963_ & ~new_n3968_;
  assign new_n3970_ = new_n3960_ & ~new_n3969_;
  assign new_n3971_ = ~new_n3960_ & new_n3969_;
  assign new_n3972_ = ~new_n3970_ & ~new_n3971_;
  assign new_n3973_ = ~new_n3486_ & ~new_n3972_;
  assign new_n3974_ = new_n3486_ & new_n3972_;
  assign new_n3975_ = ~new_n3973_ & ~new_n3974_;
  assign miter = new_n3432_ & new_n3975_;
endmodule


