// Benchmark "cir1_cir2_miter" written by ABC on Tue Jul 11 18:28:49 2023

module cir1_cir2_miter ( 
    \i:n2_control_0 , \i:n2_control_1 , \i:n2_control_2 , \i:n2_control_3 ,
    \i:n2_control_4 , \i:n4_control_0 , \i:n4_control_1 , \i:n4_control_2 ,
    \i:n4_control_3 , \i:n4_control_4 , \i:n12_control_0 ,
    \i:n12_control_1 , \i:n12_control_2 , \i:n12_control_3 ,
    \i:n12_control_4 , \i:n18_control_0 , \i:n18_control_1 ,
    \i:n18_control_2 , \i:n18_control_3 , \i:n18_control_4 ,
    \i:n22_control_0 , \i:n22_control_1 , \i:n22_control_2 ,
    \i:n22_control_3 , \i:n22_control_4 , \i:n34_control_0 ,
    \i:n34_control_1 , \i:n34_control_2 , \i:n34_control_3 ,
    \i:n34_control_4 , \i:n35_control_0 , \i:n35_control_1 ,
    \i:n35_control_2 , \i:n35_control_3 , \i:n35_control_4 ,
    \i:n51_control_0 , \i:n51_control_1 , \i:n51_control_2 ,
    \i:n51_control_3 , \i:n51_control_4 , \i:n57_control_0 ,
    \i:n57_control_1 , \i:n57_control_2 , \i:n57_control_3 ,
    \i:n57_control_4 , \i:n67_control_0 , \i:n67_control_1 ,
    \i:n67_control_2 , \i:n67_control_3 , \i:n67_control_4 ,
    \i:n72_control_0 , \i:n72_control_1 , \i:n72_control_2 ,
    \i:n72_control_3 , \i:n72_control_4 , \i:n75_control_0 ,
    \i:n75_control_1 , \i:n75_control_2 , \i:n75_control_3 ,
    \i:n75_control_4 , \i:n78_control_0 , \i:n78_control_1 ,
    \i:n78_control_2 , \i:n78_control_3 , \i:n78_control_4 ,
    \i:n80_control_0 , \i:n80_control_1 , \i:n80_control_2 ,
    \i:n80_control_3 , \i:n80_control_4 , \o:n6->n4 , \o:~n6->n4 ,
    \o:n6->n10 , \o:~n6->n10 , \o:n6->n33 , \o:~n6->n33 , \o:n6->n39 ,
    \o:~n6->n39 , \o:n6->n66 , \o:~n6->n66 , \o:n6->n70 , \o:~n6->n70 ,
    \o:n6->n71 , \o:~n6->n71 , \o:n6->n79 , \o:~n6->n79 , \o:n9->n4 ,
    \o:~n9->n4 , \o:n9->n10 , \o:~n9->n10 , \o:n9->n33 , \o:~n9->n33 ,
    \o:n9->n39 , \o:~n9->n39 , \o:n9->n66 , \o:~n9->n66 , \o:n9->n70 ,
    \o:~n9->n70 , \o:n9->n71 , \o:~n9->n71 , \o:n9->n79 , \o:~n9->n79 ,
    \o:n42->n4 , \o:~n42->n4 , \o:n42->n10 , \o:~n42->n10 , \o:n42->n33 ,
    \o:~n42->n33 , \o:n42->n39 , \o:~n42->n39 , \o:n42->n66 ,
    \o:~n42->n66 , \o:n42->n70 , \o:~n42->n70 , \o:n42->n71 ,
    \o:~n42->n71 , \o:n42->n79 , \o:~n42->n79 , \o:n48->n4 , \o:~n48->n4 ,
    \o:n48->n10 , \o:~n48->n10 , \o:n48->n33 , \o:~n48->n33 , \o:n48->n39 ,
    \o:~n48->n39 , \o:n48->n66 , \o:~n48->n66 , \o:n48->n70 ,
    \o:~n48->n70 , \o:n48->n71 , \o:~n48->n71 , \o:n48->n79 ,
    \o:~n48->n79 , \o:n56->n4 , \o:~n56->n4 , \o:n56->n10 , \o:~n56->n10 ,
    \o:n56->n33 , \o:~n56->n33 , \o:n56->n39 , \o:~n56->n39 , \o:n56->n66 ,
    \o:~n56->n66 , \o:n56->n70 , \o:~n56->n70 , \o:n56->n71 ,
    \o:~n56->n71 , \o:n56->n79 , \o:~n56->n79 , \o:n65->n4 , \o:~n65->n4 ,
    \o:n65->n10 , \o:~n65->n10 , \o:n65->n33 , \o:~n65->n33 , \o:n65->n39 ,
    \o:~n65->n39 , \o:n65->n66 , \o:~n65->n66 , \o:n65->n70 ,
    \o:~n65->n70 , \o:n65->n71 , \o:~n65->n71 , \o:n65->n79 ,
    \o:~n65->n79 , \o:n68->n4 , \o:~n68->n4 , \o:n68->n10 , \o:~n68->n10 ,
    \o:n68->n33 , \o:~n68->n33 , \o:n68->n39 , \o:~n68->n39 , \o:n68->n66 ,
    \o:~n68->n66 , \o:n68->n70 , \o:~n68->n70 , \o:n68->n71 ,
    \o:~n68->n71 , \o:n68->n79 , \o:~n68->n79 , \o:n77->n4 , \o:~n77->n4 ,
    \o:n77->n10 , \o:~n77->n10 , \o:n77->n33 , \o:~n77->n33 , \o:n77->n39 ,
    \o:~n77->n39 , \o:n77->n66 , \o:~n77->n66 , \o:n77->n70 ,
    \o:~n77->n70 , \o:n77->n71 , \o:~n77->n71 , \o:n77->n79 ,
    \o:~n77->n79 , n0_ntk1, n3_ntk1, n11_ntk1, n15_ntk1, n21_ntk1,
    n35_ntk1, n36_ntk1, n37_ntk1, n41_ntk1, n61_ntk1, n73_ntk1, n80_ntk1,
    n4381  );
  input  \i:n2_control_0 , \i:n2_control_1 , \i:n2_control_2 ,
    \i:n2_control_3 , \i:n2_control_4 , \i:n4_control_0 , \i:n4_control_1 ,
    \i:n4_control_2 , \i:n4_control_3 , \i:n4_control_4 ,
    \i:n12_control_0 , \i:n12_control_1 , \i:n12_control_2 ,
    \i:n12_control_3 , \i:n12_control_4 , \i:n18_control_0 ,
    \i:n18_control_1 , \i:n18_control_2 , \i:n18_control_3 ,
    \i:n18_control_4 , \i:n22_control_0 , \i:n22_control_1 ,
    \i:n22_control_2 , \i:n22_control_3 , \i:n22_control_4 ,
    \i:n34_control_0 , \i:n34_control_1 , \i:n34_control_2 ,
    \i:n34_control_3 , \i:n34_control_4 , \i:n35_control_0 ,
    \i:n35_control_1 , \i:n35_control_2 , \i:n35_control_3 ,
    \i:n35_control_4 , \i:n51_control_0 , \i:n51_control_1 ,
    \i:n51_control_2 , \i:n51_control_3 , \i:n51_control_4 ,
    \i:n57_control_0 , \i:n57_control_1 , \i:n57_control_2 ,
    \i:n57_control_3 , \i:n57_control_4 , \i:n67_control_0 ,
    \i:n67_control_1 , \i:n67_control_2 , \i:n67_control_3 ,
    \i:n67_control_4 , \i:n72_control_0 , \i:n72_control_1 ,
    \i:n72_control_2 , \i:n72_control_3 , \i:n72_control_4 ,
    \i:n75_control_0 , \i:n75_control_1 , \i:n75_control_2 ,
    \i:n75_control_3 , \i:n75_control_4 , \i:n78_control_0 ,
    \i:n78_control_1 , \i:n78_control_2 , \i:n78_control_3 ,
    \i:n78_control_4 , \i:n80_control_0 , \i:n80_control_1 ,
    \i:n80_control_2 , \i:n80_control_3 , \i:n80_control_4 , \o:n6->n4 ,
    \o:~n6->n4 , \o:n6->n10 , \o:~n6->n10 , \o:n6->n33 , \o:~n6->n33 ,
    \o:n6->n39 , \o:~n6->n39 , \o:n6->n66 , \o:~n6->n66 , \o:n6->n70 ,
    \o:~n6->n70 , \o:n6->n71 , \o:~n6->n71 , \o:n6->n79 , \o:~n6->n79 ,
    \o:n9->n4 , \o:~n9->n4 , \o:n9->n10 , \o:~n9->n10 , \o:n9->n33 ,
    \o:~n9->n33 , \o:n9->n39 , \o:~n9->n39 , \o:n9->n66 , \o:~n9->n66 ,
    \o:n9->n70 , \o:~n9->n70 , \o:n9->n71 , \o:~n9->n71 , \o:n9->n79 ,
    \o:~n9->n79 , \o:n42->n4 , \o:~n42->n4 , \o:n42->n10 , \o:~n42->n10 ,
    \o:n42->n33 , \o:~n42->n33 , \o:n42->n39 , \o:~n42->n39 , \o:n42->n66 ,
    \o:~n42->n66 , \o:n42->n70 , \o:~n42->n70 , \o:n42->n71 ,
    \o:~n42->n71 , \o:n42->n79 , \o:~n42->n79 , \o:n48->n4 , \o:~n48->n4 ,
    \o:n48->n10 , \o:~n48->n10 , \o:n48->n33 , \o:~n48->n33 , \o:n48->n39 ,
    \o:~n48->n39 , \o:n48->n66 , \o:~n48->n66 , \o:n48->n70 ,
    \o:~n48->n70 , \o:n48->n71 , \o:~n48->n71 , \o:n48->n79 ,
    \o:~n48->n79 , \o:n56->n4 , \o:~n56->n4 , \o:n56->n10 , \o:~n56->n10 ,
    \o:n56->n33 , \o:~n56->n33 , \o:n56->n39 , \o:~n56->n39 , \o:n56->n66 ,
    \o:~n56->n66 , \o:n56->n70 , \o:~n56->n70 , \o:n56->n71 ,
    \o:~n56->n71 , \o:n56->n79 , \o:~n56->n79 , \o:n65->n4 , \o:~n65->n4 ,
    \o:n65->n10 , \o:~n65->n10 , \o:n65->n33 , \o:~n65->n33 , \o:n65->n39 ,
    \o:~n65->n39 , \o:n65->n66 , \o:~n65->n66 , \o:n65->n70 ,
    \o:~n65->n70 , \o:n65->n71 , \o:~n65->n71 , \o:n65->n79 ,
    \o:~n65->n79 , \o:n68->n4 , \o:~n68->n4 , \o:n68->n10 , \o:~n68->n10 ,
    \o:n68->n33 , \o:~n68->n33 , \o:n68->n39 , \o:~n68->n39 , \o:n68->n66 ,
    \o:~n68->n66 , \o:n68->n70 , \o:~n68->n70 , \o:n68->n71 ,
    \o:~n68->n71 , \o:n68->n79 , \o:~n68->n79 , \o:n77->n4 , \o:~n77->n4 ,
    \o:n77->n10 , \o:~n77->n10 , \o:n77->n33 , \o:~n77->n33 , \o:n77->n39 ,
    \o:~n77->n39 , \o:n77->n66 , \o:~n77->n66 , \o:n77->n70 ,
    \o:~n77->n70 , \o:n77->n71 , \o:~n77->n71 , \o:n77->n79 ,
    \o:~n77->n79 , n0_ntk1, n3_ntk1, n11_ntk1, n15_ntk1, n21_ntk1,
    n35_ntk1, n36_ntk1, n37_ntk1, n41_ntk1, n61_ntk1, n73_ntk1, n80_ntk1;
  output n4381;
  wire new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_,
    new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_,
    new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_,
    new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_,
    new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_,
    new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_,
    new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_,
    new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_,
    new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_,
    new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_,
    new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_,
    new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_,
    new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_,
    new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_,
    new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_,
    new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_,
    new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_,
    new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_,
    new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_,
    new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_,
    new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_,
    new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_,
    new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_,
    new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_,
    new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_,
    new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_,
    new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_,
    new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_,
    new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_,
    new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_,
    new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_,
    new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_,
    new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_,
    new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_,
    new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_,
    new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_,
    new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_,
    new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_,
    new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_,
    new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_,
    new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_,
    new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_,
    new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_,
    new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_,
    new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_,
    new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_,
    new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_,
    new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_,
    new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_,
    new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_,
    new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_,
    new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_,
    new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_,
    new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_,
    new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_,
    new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_,
    new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_,
    new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_,
    new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_,
    new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_,
    new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_,
    new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_,
    new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_,
    new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_,
    new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_,
    new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_,
    new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_,
    new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_,
    new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_,
    new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_,
    new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_,
    new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_,
    new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_,
    new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_,
    new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_,
    new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_,
    new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_,
    new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_,
    new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_,
    new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_,
    new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_,
    new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_,
    new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_,
    new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_,
    new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_,
    new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_,
    new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_,
    new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_,
    new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_,
    new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_,
    new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_,
    new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_,
    new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_,
    new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_,
    new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_,
    new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_,
    new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_,
    new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_,
    new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_,
    new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_,
    new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_,
    new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_,
    new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_,
    new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_,
    new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_,
    new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_,
    new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_,
    new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_,
    new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_,
    new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_,
    new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_,
    new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_,
    new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_,
    new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_,
    new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_,
    new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_,
    new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_,
    new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_,
    new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_,
    new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_,
    new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_,
    new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_,
    new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_,
    new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_,
    new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_,
    new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_,
    new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_,
    new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_,
    new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_,
    new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_,
    new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_,
    new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_,
    new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_,
    new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_,
    new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_,
    new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_,
    new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_,
    new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_,
    new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_,
    new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_,
    new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_,
    new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_,
    new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_,
    new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_,
    new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_,
    new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_,
    new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1741_,
    new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_,
    new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_,
    new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_, new_n1759_,
    new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_, new_n1765_,
    new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_,
    new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1777_,
    new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_, new_n1783_,
    new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_,
    new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_,
    new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_,
    new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_,
    new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_,
    new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_,
    new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_,
    new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_,
    new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_,
    new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_,
    new_n1844_, new_n1845_;
  assign new_n212_ = n3_ntk1 & ~n80_ntk1;
  assign new_n213_ = ~n3_ntk1 & ~n41_ntk1;
  assign new_n214_ = ~new_n212_ & ~new_n213_;
  assign new_n215_ = ~n37_ntk1 & ~new_n214_;
  assign new_n216_ = ~n3_ntk1 & n21_ntk1;
  assign new_n217_ = n3_ntk1 & n73_ntk1;
  assign new_n218_ = ~new_n216_ & ~new_n217_;
  assign new_n219_ = n37_ntk1 & ~new_n218_;
  assign new_n220_ = n21_ntk1 & ~n61_ntk1;
  assign new_n221_ = n61_ntk1 & n73_ntk1;
  assign new_n222_ = ~new_n220_ & ~new_n221_;
  assign new_n223_ = n36_ntk1 & ~new_n222_;
  assign new_n224_ = ~new_n219_ & ~new_n223_;
  assign new_n225_ = ~n0_ntk1 & ~n41_ntk1;
  assign new_n226_ = n0_ntk1 & ~n80_ntk1;
  assign new_n227_ = ~new_n225_ & ~new_n226_;
  assign new_n228_ = ~n15_ntk1 & ~new_n227_;
  assign new_n229_ = ~n0_ntk1 & n21_ntk1;
  assign new_n230_ = n0_ntk1 & n73_ntk1;
  assign new_n231_ = ~new_n229_ & ~new_n230_;
  assign new_n232_ = n15_ntk1 & ~new_n231_;
  assign new_n233_ = ~n35_ntk1 & ~n41_ntk1;
  assign new_n234_ = n35_ntk1 & ~n80_ntk1;
  assign new_n235_ = ~new_n233_ & ~new_n234_;
  assign new_n236_ = ~n11_ntk1 & ~new_n235_;
  assign new_n237_ = ~new_n232_ & new_n236_;
  assign new_n238_ = ~new_n228_ & ~new_n237_;
  assign new_n239_ = new_n224_ & ~new_n238_;
  assign new_n240_ = ~n41_ntk1 & ~n61_ntk1;
  assign new_n241_ = n61_ntk1 & ~n80_ntk1;
  assign new_n242_ = ~new_n240_ & ~new_n241_;
  assign new_n243_ = ~n36_ntk1 & ~new_n242_;
  assign new_n244_ = ~new_n219_ & new_n243_;
  assign new_n245_ = ~new_n239_ & ~new_n244_;
  assign new_n246_ = ~new_n215_ & new_n245_;
  assign new_n247_ = \i:n35_control_1  & n61_ntk1;
  assign new_n248_ = ~\i:n35_control_1  & n41_ntk1;
  assign new_n249_ = ~new_n247_ & ~new_n248_;
  assign new_n250_ = ~\i:n35_control_2  & new_n249_;
  assign new_n251_ = \i:n35_control_1  & n80_ntk1;
  assign new_n252_ = ~\i:n35_control_1  & n73_ntk1;
  assign new_n253_ = ~new_n251_ & ~new_n252_;
  assign new_n254_ = \i:n35_control_2  & new_n253_;
  assign new_n255_ = ~new_n250_ & ~new_n254_;
  assign new_n256_ = \i:n35_control_4  & ~new_n255_;
  assign new_n257_ = \i:n35_control_1  & n3_ntk1;
  assign new_n258_ = ~\i:n35_control_1  & n0_ntk1;
  assign new_n259_ = ~new_n257_ & ~new_n258_;
  assign new_n260_ = ~\i:n35_control_2  & new_n259_;
  assign new_n261_ = \i:n35_control_1  & n15_ntk1;
  assign new_n262_ = ~\i:n35_control_1  & n11_ntk1;
  assign new_n263_ = ~new_n261_ & ~new_n262_;
  assign new_n264_ = \i:n35_control_2  & new_n263_;
  assign new_n265_ = ~new_n260_ & ~new_n264_;
  assign new_n266_ = ~\i:n35_control_4  & ~new_n265_;
  assign new_n267_ = ~new_n256_ & ~new_n266_;
  assign new_n268_ = ~\i:n35_control_3  & ~new_n267_;
  assign new_n269_ = \i:n35_control_1  & n37_ntk1;
  assign new_n270_ = ~\i:n35_control_1  & n36_ntk1;
  assign new_n271_ = ~new_n269_ & ~new_n270_;
  assign new_n272_ = \i:n35_control_2  & new_n271_;
  assign new_n273_ = \i:n35_control_1  & n35_ntk1;
  assign new_n274_ = ~\i:n35_control_1  & n21_ntk1;
  assign new_n275_ = ~new_n273_ & ~new_n274_;
  assign new_n276_ = ~\i:n35_control_2  & new_n275_;
  assign new_n277_ = ~new_n272_ & ~new_n276_;
  assign new_n278_ = \i:n35_control_3  & ~new_n277_;
  assign new_n279_ = ~\i:n35_control_4  & new_n278_;
  assign new_n280_ = ~new_n268_ & ~new_n279_;
  assign new_n281_ = \i:n35_control_0  & ~new_n280_;
  assign new_n282_ = ~\i:n35_control_0  & new_n280_;
  assign new_n283_ = ~new_n281_ & ~new_n282_;
  assign new_n284_ = \i:n4_control_1  & n61_ntk1;
  assign new_n285_ = ~\i:n4_control_1  & n41_ntk1;
  assign new_n286_ = ~new_n284_ & ~new_n285_;
  assign new_n287_ = ~\i:n4_control_2  & new_n286_;
  assign new_n288_ = \i:n4_control_1  & n80_ntk1;
  assign new_n289_ = ~\i:n4_control_1  & n73_ntk1;
  assign new_n290_ = ~new_n288_ & ~new_n289_;
  assign new_n291_ = \i:n4_control_2  & new_n290_;
  assign new_n292_ = ~new_n287_ & ~new_n291_;
  assign new_n293_ = \i:n4_control_4  & ~new_n292_;
  assign new_n294_ = \i:n4_control_1  & n3_ntk1;
  assign new_n295_ = ~\i:n4_control_1  & n0_ntk1;
  assign new_n296_ = ~new_n294_ & ~new_n295_;
  assign new_n297_ = ~\i:n4_control_2  & new_n296_;
  assign new_n298_ = \i:n4_control_1  & n15_ntk1;
  assign new_n299_ = ~\i:n4_control_1  & n11_ntk1;
  assign new_n300_ = ~new_n298_ & ~new_n299_;
  assign new_n301_ = \i:n4_control_2  & new_n300_;
  assign new_n302_ = ~new_n297_ & ~new_n301_;
  assign new_n303_ = ~\i:n4_control_4  & ~new_n302_;
  assign new_n304_ = ~new_n293_ & ~new_n303_;
  assign new_n305_ = ~\i:n4_control_3  & ~new_n304_;
  assign new_n306_ = \i:n4_control_1  & n37_ntk1;
  assign new_n307_ = ~\i:n4_control_1  & n36_ntk1;
  assign new_n308_ = ~new_n306_ & ~new_n307_;
  assign new_n309_ = \i:n4_control_2  & new_n308_;
  assign new_n310_ = \i:n4_control_1  & n35_ntk1;
  assign new_n311_ = ~\i:n4_control_1  & n21_ntk1;
  assign new_n312_ = ~new_n310_ & ~new_n311_;
  assign new_n313_ = ~\i:n4_control_2  & new_n312_;
  assign new_n314_ = ~new_n309_ & ~new_n313_;
  assign new_n315_ = \i:n4_control_3  & ~new_n314_;
  assign new_n316_ = ~\i:n4_control_4  & new_n315_;
  assign new_n317_ = ~new_n305_ & ~new_n316_;
  assign new_n318_ = \i:n4_control_0  & ~new_n317_;
  assign new_n319_ = ~\i:n4_control_0  & new_n317_;
  assign new_n320_ = ~new_n318_ & ~new_n319_;
  assign new_n321_ = ~\i:n72_control_1  & ~n73_ntk1;
  assign new_n322_ = \i:n72_control_1  & ~n80_ntk1;
  assign new_n323_ = ~new_n321_ & ~new_n322_;
  assign new_n324_ = \i:n72_control_2  & ~new_n323_;
  assign new_n325_ = ~\i:n72_control_1  & ~n35_ntk1;
  assign new_n326_ = \i:n72_control_1  & ~n41_ntk1;
  assign new_n327_ = ~new_n325_ & ~new_n326_;
  assign new_n328_ = ~\i:n72_control_2  & ~new_n327_;
  assign new_n329_ = ~new_n324_ & ~new_n328_;
  assign new_n330_ = \i:n72_control_3  & ~new_n329_;
  assign new_n331_ = ~\i:n72_control_1  & ~n15_ntk1;
  assign new_n332_ = \i:n72_control_1  & ~n21_ntk1;
  assign new_n333_ = ~new_n331_ & ~new_n332_;
  assign new_n334_ = \i:n72_control_2  & ~new_n333_;
  assign new_n335_ = ~\i:n72_control_1  & ~n0_ntk1;
  assign new_n336_ = \i:n72_control_1  & ~n11_ntk1;
  assign new_n337_ = ~new_n335_ & ~new_n336_;
  assign new_n338_ = ~\i:n72_control_2  & ~new_n337_;
  assign new_n339_ = ~new_n334_ & ~new_n338_;
  assign new_n340_ = ~\i:n72_control_3  & ~new_n339_;
  assign new_n341_ = ~new_n330_ & ~new_n340_;
  assign new_n342_ = ~\i:n72_control_4  & ~new_n341_;
  assign new_n343_ = \i:n72_control_0  & new_n342_;
  assign new_n344_ = ~\i:n72_control_0  & ~new_n342_;
  assign new_n345_ = ~new_n343_ & ~new_n344_;
  assign new_n346_ = ~new_n320_ & new_n345_;
  assign new_n347_ = ~\i:n75_control_1  & ~n73_ntk1;
  assign new_n348_ = \i:n75_control_1  & ~n80_ntk1;
  assign new_n349_ = ~new_n347_ & ~new_n348_;
  assign new_n350_ = \i:n75_control_2  & ~new_n349_;
  assign new_n351_ = ~\i:n75_control_1  & ~n35_ntk1;
  assign new_n352_ = \i:n75_control_1  & ~n41_ntk1;
  assign new_n353_ = ~new_n351_ & ~new_n352_;
  assign new_n354_ = ~\i:n75_control_2  & ~new_n353_;
  assign new_n355_ = ~new_n350_ & ~new_n354_;
  assign new_n356_ = \i:n75_control_3  & ~new_n355_;
  assign new_n357_ = ~\i:n75_control_1  & ~n15_ntk1;
  assign new_n358_ = \i:n75_control_1  & ~n21_ntk1;
  assign new_n359_ = ~new_n357_ & ~new_n358_;
  assign new_n360_ = \i:n75_control_2  & ~new_n359_;
  assign new_n361_ = ~\i:n75_control_1  & ~n0_ntk1;
  assign new_n362_ = \i:n75_control_1  & ~n11_ntk1;
  assign new_n363_ = ~new_n361_ & ~new_n362_;
  assign new_n364_ = ~\i:n75_control_2  & ~new_n363_;
  assign new_n365_ = ~new_n360_ & ~new_n364_;
  assign new_n366_ = ~\i:n75_control_3  & ~new_n365_;
  assign new_n367_ = ~new_n356_ & ~new_n366_;
  assign new_n368_ = ~\i:n75_control_4  & ~new_n367_;
  assign new_n369_ = \i:n75_control_0  & new_n368_;
  assign new_n370_ = ~\i:n75_control_0  & ~new_n368_;
  assign new_n371_ = ~new_n369_ & ~new_n370_;
  assign new_n372_ = new_n320_ & new_n371_;
  assign new_n373_ = ~new_n346_ & ~new_n372_;
  assign new_n374_ = new_n283_ & ~new_n373_;
  assign new_n375_ = ~\i:n78_control_1  & ~n73_ntk1;
  assign new_n376_ = \i:n78_control_1  & ~n80_ntk1;
  assign new_n377_ = ~new_n375_ & ~new_n376_;
  assign new_n378_ = \i:n78_control_2  & ~new_n377_;
  assign new_n379_ = ~\i:n78_control_1  & ~n35_ntk1;
  assign new_n380_ = \i:n78_control_1  & ~n41_ntk1;
  assign new_n381_ = ~new_n379_ & ~new_n380_;
  assign new_n382_ = ~\i:n78_control_2  & ~new_n381_;
  assign new_n383_ = ~new_n378_ & ~new_n382_;
  assign new_n384_ = \i:n78_control_3  & ~new_n383_;
  assign new_n385_ = ~\i:n78_control_1  & ~n15_ntk1;
  assign new_n386_ = \i:n78_control_1  & ~n21_ntk1;
  assign new_n387_ = ~new_n385_ & ~new_n386_;
  assign new_n388_ = \i:n78_control_2  & ~new_n387_;
  assign new_n389_ = ~\i:n78_control_1  & ~n0_ntk1;
  assign new_n390_ = \i:n78_control_1  & ~n11_ntk1;
  assign new_n391_ = ~new_n389_ & ~new_n390_;
  assign new_n392_ = ~\i:n78_control_2  & ~new_n391_;
  assign new_n393_ = ~new_n388_ & ~new_n392_;
  assign new_n394_ = ~\i:n78_control_3  & ~new_n393_;
  assign new_n395_ = ~new_n384_ & ~new_n394_;
  assign new_n396_ = ~\i:n78_control_4  & ~new_n395_;
  assign new_n397_ = \i:n78_control_0  & new_n396_;
  assign new_n398_ = ~\i:n78_control_0  & ~new_n396_;
  assign new_n399_ = ~new_n397_ & ~new_n398_;
  assign new_n400_ = ~new_n320_ & ~new_n399_;
  assign new_n401_ = ~\i:n80_control_1  & ~n73_ntk1;
  assign new_n402_ = \i:n80_control_1  & ~n80_ntk1;
  assign new_n403_ = ~new_n401_ & ~new_n402_;
  assign new_n404_ = \i:n80_control_2  & ~new_n403_;
  assign new_n405_ = ~\i:n80_control_1  & ~n35_ntk1;
  assign new_n406_ = \i:n80_control_1  & ~n41_ntk1;
  assign new_n407_ = ~new_n405_ & ~new_n406_;
  assign new_n408_ = ~\i:n80_control_2  & ~new_n407_;
  assign new_n409_ = ~new_n404_ & ~new_n408_;
  assign new_n410_ = \i:n80_control_3  & ~new_n409_;
  assign new_n411_ = ~\i:n80_control_1  & ~n15_ntk1;
  assign new_n412_ = \i:n80_control_1  & ~n21_ntk1;
  assign new_n413_ = ~new_n411_ & ~new_n412_;
  assign new_n414_ = \i:n80_control_2  & ~new_n413_;
  assign new_n415_ = ~\i:n80_control_1  & ~n0_ntk1;
  assign new_n416_ = \i:n80_control_1  & ~n11_ntk1;
  assign new_n417_ = ~new_n415_ & ~new_n416_;
  assign new_n418_ = ~\i:n80_control_2  & ~new_n417_;
  assign new_n419_ = ~new_n414_ & ~new_n418_;
  assign new_n420_ = ~\i:n80_control_3  & ~new_n419_;
  assign new_n421_ = ~new_n410_ & ~new_n420_;
  assign new_n422_ = ~\i:n80_control_4  & ~new_n421_;
  assign new_n423_ = \i:n80_control_0  & new_n422_;
  assign new_n424_ = ~\i:n80_control_0  & ~new_n422_;
  assign new_n425_ = ~new_n423_ & ~new_n424_;
  assign new_n426_ = new_n320_ & ~new_n425_;
  assign new_n427_ = ~new_n400_ & ~new_n426_;
  assign new_n428_ = ~new_n283_ & ~new_n427_;
  assign new_n429_ = \i:n34_control_1  & n61_ntk1;
  assign new_n430_ = ~\i:n34_control_1  & n41_ntk1;
  assign new_n431_ = ~new_n429_ & ~new_n430_;
  assign new_n432_ = ~\i:n34_control_2  & new_n431_;
  assign new_n433_ = \i:n34_control_1  & n80_ntk1;
  assign new_n434_ = ~\i:n34_control_1  & n73_ntk1;
  assign new_n435_ = ~new_n433_ & ~new_n434_;
  assign new_n436_ = \i:n34_control_2  & new_n435_;
  assign new_n437_ = ~new_n432_ & ~new_n436_;
  assign new_n438_ = \i:n34_control_4  & ~new_n437_;
  assign new_n439_ = \i:n34_control_1  & n3_ntk1;
  assign new_n440_ = ~\i:n34_control_1  & n0_ntk1;
  assign new_n441_ = ~new_n439_ & ~new_n440_;
  assign new_n442_ = ~\i:n34_control_2  & new_n441_;
  assign new_n443_ = \i:n34_control_1  & n15_ntk1;
  assign new_n444_ = ~\i:n34_control_1  & n11_ntk1;
  assign new_n445_ = ~new_n443_ & ~new_n444_;
  assign new_n446_ = \i:n34_control_2  & new_n445_;
  assign new_n447_ = ~new_n442_ & ~new_n446_;
  assign new_n448_ = ~\i:n34_control_4  & ~new_n447_;
  assign new_n449_ = ~new_n438_ & ~new_n448_;
  assign new_n450_ = ~\i:n34_control_3  & ~new_n449_;
  assign new_n451_ = \i:n34_control_1  & n37_ntk1;
  assign new_n452_ = ~\i:n34_control_1  & n36_ntk1;
  assign new_n453_ = ~new_n451_ & ~new_n452_;
  assign new_n454_ = \i:n34_control_2  & new_n453_;
  assign new_n455_ = \i:n34_control_1  & n35_ntk1;
  assign new_n456_ = ~\i:n34_control_1  & n21_ntk1;
  assign new_n457_ = ~new_n455_ & ~new_n456_;
  assign new_n458_ = ~\i:n34_control_2  & new_n457_;
  assign new_n459_ = ~new_n454_ & ~new_n458_;
  assign new_n460_ = \i:n34_control_3  & ~new_n459_;
  assign new_n461_ = ~\i:n34_control_4  & new_n460_;
  assign new_n462_ = ~new_n450_ & ~new_n461_;
  assign new_n463_ = \i:n34_control_0  & ~new_n462_;
  assign new_n464_ = ~\i:n34_control_0  & new_n462_;
  assign new_n465_ = ~new_n463_ & ~new_n464_;
  assign new_n466_ = \i:n57_control_1  & n61_ntk1;
  assign new_n467_ = ~\i:n57_control_1  & n41_ntk1;
  assign new_n468_ = ~new_n466_ & ~new_n467_;
  assign new_n469_ = ~\i:n57_control_2  & new_n468_;
  assign new_n470_ = \i:n57_control_1  & n80_ntk1;
  assign new_n471_ = ~\i:n57_control_1  & n73_ntk1;
  assign new_n472_ = ~new_n470_ & ~new_n471_;
  assign new_n473_ = \i:n57_control_2  & new_n472_;
  assign new_n474_ = ~new_n469_ & ~new_n473_;
  assign new_n475_ = \i:n57_control_4  & ~new_n474_;
  assign new_n476_ = \i:n57_control_1  & n3_ntk1;
  assign new_n477_ = ~\i:n57_control_1  & n0_ntk1;
  assign new_n478_ = ~new_n476_ & ~new_n477_;
  assign new_n479_ = ~\i:n57_control_2  & new_n478_;
  assign new_n480_ = \i:n57_control_1  & n15_ntk1;
  assign new_n481_ = ~\i:n57_control_1  & n11_ntk1;
  assign new_n482_ = ~new_n480_ & ~new_n481_;
  assign new_n483_ = \i:n57_control_2  & new_n482_;
  assign new_n484_ = ~new_n479_ & ~new_n483_;
  assign new_n485_ = ~\i:n57_control_4  & ~new_n484_;
  assign new_n486_ = ~new_n475_ & ~new_n485_;
  assign new_n487_ = ~\i:n57_control_3  & ~new_n486_;
  assign new_n488_ = \i:n57_control_1  & n37_ntk1;
  assign new_n489_ = ~\i:n57_control_1  & n36_ntk1;
  assign new_n490_ = ~new_n488_ & ~new_n489_;
  assign new_n491_ = \i:n57_control_2  & new_n490_;
  assign new_n492_ = \i:n57_control_1  & n35_ntk1;
  assign new_n493_ = ~\i:n57_control_1  & n21_ntk1;
  assign new_n494_ = ~new_n492_ & ~new_n493_;
  assign new_n495_ = ~\i:n57_control_2  & new_n494_;
  assign new_n496_ = ~new_n491_ & ~new_n495_;
  assign new_n497_ = \i:n57_control_3  & ~new_n496_;
  assign new_n498_ = ~\i:n57_control_4  & new_n497_;
  assign new_n499_ = ~new_n487_ & ~new_n498_;
  assign new_n500_ = \i:n57_control_0  & ~new_n499_;
  assign new_n501_ = ~\i:n57_control_0  & new_n499_;
  assign new_n502_ = ~new_n500_ & ~new_n501_;
  assign new_n503_ = new_n345_ & ~new_n502_;
  assign new_n504_ = new_n371_ & new_n502_;
  assign new_n505_ = ~new_n503_ & ~new_n504_;
  assign new_n506_ = new_n465_ & ~new_n505_;
  assign new_n507_ = \i:n18_control_1  & n61_ntk1;
  assign new_n508_ = ~\i:n18_control_1  & n41_ntk1;
  assign new_n509_ = ~new_n507_ & ~new_n508_;
  assign new_n510_ = ~\i:n18_control_2  & new_n509_;
  assign new_n511_ = \i:n18_control_1  & n80_ntk1;
  assign new_n512_ = ~\i:n18_control_1  & n73_ntk1;
  assign new_n513_ = ~new_n511_ & ~new_n512_;
  assign new_n514_ = \i:n18_control_2  & new_n513_;
  assign new_n515_ = ~new_n510_ & ~new_n514_;
  assign new_n516_ = \i:n18_control_4  & ~new_n515_;
  assign new_n517_ = \i:n18_control_1  & n3_ntk1;
  assign new_n518_ = ~\i:n18_control_1  & n0_ntk1;
  assign new_n519_ = ~new_n517_ & ~new_n518_;
  assign new_n520_ = ~\i:n18_control_2  & new_n519_;
  assign new_n521_ = \i:n18_control_1  & n15_ntk1;
  assign new_n522_ = ~\i:n18_control_1  & n11_ntk1;
  assign new_n523_ = ~new_n521_ & ~new_n522_;
  assign new_n524_ = \i:n18_control_2  & new_n523_;
  assign new_n525_ = ~new_n520_ & ~new_n524_;
  assign new_n526_ = ~\i:n18_control_4  & ~new_n525_;
  assign new_n527_ = ~new_n516_ & ~new_n526_;
  assign new_n528_ = ~\i:n18_control_3  & ~new_n527_;
  assign new_n529_ = \i:n18_control_1  & n37_ntk1;
  assign new_n530_ = ~\i:n18_control_1  & n36_ntk1;
  assign new_n531_ = ~new_n529_ & ~new_n530_;
  assign new_n532_ = \i:n18_control_2  & new_n531_;
  assign new_n533_ = \i:n18_control_1  & n35_ntk1;
  assign new_n534_ = ~\i:n18_control_1  & n21_ntk1;
  assign new_n535_ = ~new_n533_ & ~new_n534_;
  assign new_n536_ = ~\i:n18_control_2  & new_n535_;
  assign new_n537_ = ~new_n532_ & ~new_n536_;
  assign new_n538_ = \i:n18_control_3  & ~new_n537_;
  assign new_n539_ = ~\i:n18_control_4  & new_n538_;
  assign new_n540_ = ~new_n528_ & ~new_n539_;
  assign new_n541_ = \i:n18_control_0  & ~new_n540_;
  assign new_n542_ = ~\i:n18_control_0  & new_n540_;
  assign new_n543_ = ~new_n541_ & ~new_n542_;
  assign new_n544_ = \i:n2_control_1  & n61_ntk1;
  assign new_n545_ = ~\i:n2_control_1  & n41_ntk1;
  assign new_n546_ = ~new_n544_ & ~new_n545_;
  assign new_n547_ = ~\i:n2_control_2  & new_n546_;
  assign new_n548_ = \i:n2_control_1  & n80_ntk1;
  assign new_n549_ = ~\i:n2_control_1  & n73_ntk1;
  assign new_n550_ = ~new_n548_ & ~new_n549_;
  assign new_n551_ = \i:n2_control_2  & new_n550_;
  assign new_n552_ = ~new_n547_ & ~new_n551_;
  assign new_n553_ = \i:n2_control_4  & ~new_n552_;
  assign new_n554_ = \i:n2_control_1  & n3_ntk1;
  assign new_n555_ = ~\i:n2_control_1  & n0_ntk1;
  assign new_n556_ = ~new_n554_ & ~new_n555_;
  assign new_n557_ = ~\i:n2_control_2  & new_n556_;
  assign new_n558_ = \i:n2_control_1  & n15_ntk1;
  assign new_n559_ = ~\i:n2_control_1  & n11_ntk1;
  assign new_n560_ = ~new_n558_ & ~new_n559_;
  assign new_n561_ = \i:n2_control_2  & new_n560_;
  assign new_n562_ = ~new_n557_ & ~new_n561_;
  assign new_n563_ = ~\i:n2_control_4  & ~new_n562_;
  assign new_n564_ = ~new_n553_ & ~new_n563_;
  assign new_n565_ = ~\i:n2_control_3  & ~new_n564_;
  assign new_n566_ = \i:n2_control_1  & n37_ntk1;
  assign new_n567_ = ~\i:n2_control_1  & n36_ntk1;
  assign new_n568_ = ~new_n566_ & ~new_n567_;
  assign new_n569_ = \i:n2_control_2  & new_n568_;
  assign new_n570_ = \i:n2_control_1  & n35_ntk1;
  assign new_n571_ = ~\i:n2_control_1  & n21_ntk1;
  assign new_n572_ = ~new_n570_ & ~new_n571_;
  assign new_n573_ = ~\i:n2_control_2  & new_n572_;
  assign new_n574_ = ~new_n569_ & ~new_n573_;
  assign new_n575_ = \i:n2_control_3  & ~new_n574_;
  assign new_n576_ = ~\i:n2_control_4  & new_n575_;
  assign new_n577_ = ~new_n565_ & ~new_n576_;
  assign new_n578_ = \i:n2_control_0  & ~new_n577_;
  assign new_n579_ = ~\i:n2_control_0  & new_n577_;
  assign new_n580_ = ~new_n578_ & ~new_n579_;
  assign new_n581_ = new_n345_ & ~new_n580_;
  assign new_n582_ = new_n371_ & new_n580_;
  assign new_n583_ = ~new_n581_ & ~new_n582_;
  assign new_n584_ = new_n543_ & ~new_n583_;
  assign new_n585_ = ~\i:n22_control_1  & ~n73_ntk1;
  assign new_n586_ = \i:n22_control_1  & ~n80_ntk1;
  assign new_n587_ = ~new_n585_ & ~new_n586_;
  assign new_n588_ = \i:n22_control_2  & ~new_n587_;
  assign new_n589_ = ~\i:n22_control_1  & ~n35_ntk1;
  assign new_n590_ = \i:n22_control_1  & ~n41_ntk1;
  assign new_n591_ = ~new_n589_ & ~new_n590_;
  assign new_n592_ = ~\i:n22_control_2  & ~new_n591_;
  assign new_n593_ = ~new_n588_ & ~new_n592_;
  assign new_n594_ = \i:n22_control_3  & ~new_n593_;
  assign new_n595_ = ~\i:n22_control_1  & ~n15_ntk1;
  assign new_n596_ = \i:n22_control_1  & ~n21_ntk1;
  assign new_n597_ = ~new_n595_ & ~new_n596_;
  assign new_n598_ = \i:n22_control_2  & ~new_n597_;
  assign new_n599_ = ~\i:n22_control_1  & ~n0_ntk1;
  assign new_n600_ = \i:n22_control_1  & ~n11_ntk1;
  assign new_n601_ = ~new_n599_ & ~new_n600_;
  assign new_n602_ = ~\i:n22_control_2  & ~new_n601_;
  assign new_n603_ = ~new_n598_ & ~new_n602_;
  assign new_n604_ = ~\i:n22_control_3  & ~new_n603_;
  assign new_n605_ = ~new_n594_ & ~new_n604_;
  assign new_n606_ = ~\i:n22_control_4  & ~new_n605_;
  assign new_n607_ = \i:n22_control_0  & new_n606_;
  assign new_n608_ = ~\i:n22_control_0  & ~new_n606_;
  assign new_n609_ = ~new_n607_ & ~new_n608_;
  assign new_n610_ = ~\i:n67_control_1  & ~n73_ntk1;
  assign new_n611_ = \i:n67_control_1  & ~n80_ntk1;
  assign new_n612_ = ~new_n610_ & ~new_n611_;
  assign new_n613_ = \i:n67_control_2  & ~new_n612_;
  assign new_n614_ = ~\i:n67_control_1  & ~n35_ntk1;
  assign new_n615_ = \i:n67_control_1  & ~n41_ntk1;
  assign new_n616_ = ~new_n614_ & ~new_n615_;
  assign new_n617_ = ~\i:n67_control_2  & ~new_n616_;
  assign new_n618_ = ~new_n613_ & ~new_n617_;
  assign new_n619_ = \i:n67_control_3  & ~new_n618_;
  assign new_n620_ = ~\i:n67_control_1  & ~n15_ntk1;
  assign new_n621_ = \i:n67_control_1  & ~n21_ntk1;
  assign new_n622_ = ~new_n620_ & ~new_n621_;
  assign new_n623_ = \i:n67_control_2  & ~new_n622_;
  assign new_n624_ = ~\i:n67_control_1  & ~n0_ntk1;
  assign new_n625_ = \i:n67_control_1  & ~n11_ntk1;
  assign new_n626_ = ~new_n624_ & ~new_n625_;
  assign new_n627_ = ~\i:n67_control_2  & ~new_n626_;
  assign new_n628_ = ~new_n623_ & ~new_n627_;
  assign new_n629_ = ~\i:n67_control_3  & ~new_n628_;
  assign new_n630_ = ~new_n619_ & ~new_n629_;
  assign new_n631_ = ~\i:n67_control_4  & ~new_n630_;
  assign new_n632_ = \i:n67_control_0  & new_n631_;
  assign new_n633_ = ~\i:n67_control_0  & ~new_n631_;
  assign new_n634_ = ~new_n632_ & ~new_n633_;
  assign new_n635_ = new_n345_ & ~new_n634_;
  assign new_n636_ = new_n371_ & new_n634_;
  assign new_n637_ = ~new_n635_ & ~new_n636_;
  assign new_n638_ = new_n609_ & ~new_n637_;
  assign new_n639_ = ~new_n399_ & ~new_n580_;
  assign new_n640_ = ~new_n425_ & new_n580_;
  assign new_n641_ = ~new_n639_ & ~new_n640_;
  assign new_n642_ = ~new_n543_ & ~new_n641_;
  assign new_n643_ = new_n638_ & ~new_n642_;
  assign new_n644_ = ~new_n584_ & ~new_n643_;
  assign new_n645_ = ~new_n399_ & ~new_n502_;
  assign new_n646_ = ~new_n425_ & new_n502_;
  assign new_n647_ = ~new_n645_ & ~new_n646_;
  assign new_n648_ = ~new_n465_ & ~new_n647_;
  assign new_n649_ = ~new_n644_ & ~new_n648_;
  assign new_n650_ = ~new_n506_ & ~new_n649_;
  assign new_n651_ = ~new_n428_ & ~new_n650_;
  assign new_n652_ = ~new_n374_ & ~new_n651_;
  assign new_n653_ = ~\i:n51_control_1  & ~n73_ntk1;
  assign new_n654_ = \i:n51_control_1  & ~n80_ntk1;
  assign new_n655_ = ~new_n653_ & ~new_n654_;
  assign new_n656_ = \i:n51_control_2  & ~new_n655_;
  assign new_n657_ = ~\i:n51_control_1  & ~n35_ntk1;
  assign new_n658_ = \i:n51_control_1  & ~n41_ntk1;
  assign new_n659_ = ~new_n657_ & ~new_n658_;
  assign new_n660_ = ~\i:n51_control_2  & ~new_n659_;
  assign new_n661_ = ~new_n656_ & ~new_n660_;
  assign new_n662_ = \i:n51_control_3  & ~new_n661_;
  assign new_n663_ = ~\i:n51_control_1  & ~n15_ntk1;
  assign new_n664_ = \i:n51_control_1  & ~n21_ntk1;
  assign new_n665_ = ~new_n663_ & ~new_n664_;
  assign new_n666_ = \i:n51_control_2  & ~new_n665_;
  assign new_n667_ = ~\i:n51_control_1  & ~n0_ntk1;
  assign new_n668_ = \i:n51_control_1  & ~n11_ntk1;
  assign new_n669_ = ~new_n667_ & ~new_n668_;
  assign new_n670_ = ~\i:n51_control_2  & ~new_n669_;
  assign new_n671_ = ~new_n666_ & ~new_n670_;
  assign new_n672_ = ~\i:n51_control_3  & ~new_n671_;
  assign new_n673_ = ~new_n662_ & ~new_n672_;
  assign new_n674_ = ~\i:n51_control_4  & ~new_n673_;
  assign new_n675_ = \i:n51_control_0  & new_n674_;
  assign new_n676_ = ~\i:n51_control_0  & ~new_n674_;
  assign new_n677_ = ~new_n675_ & ~new_n676_;
  assign new_n678_ = ~new_n399_ & ~new_n634_;
  assign new_n679_ = ~new_n425_ & new_n634_;
  assign new_n680_ = ~new_n678_ & ~new_n679_;
  assign new_n681_ = ~new_n609_ & ~new_n680_;
  assign new_n682_ = ~new_n642_ & ~new_n681_;
  assign new_n683_ = ~new_n428_ & ~new_n648_;
  assign new_n684_ = new_n682_ & new_n683_;
  assign new_n685_ = ~new_n677_ & new_n684_;
  assign new_n686_ = new_n652_ & ~new_n685_;
  assign new_n687_ = ~new_n246_ & new_n686_;
  assign new_n688_ = n21_ntk1 & ~n35_ntk1;
  assign new_n689_ = n35_ntk1 & n73_ntk1;
  assign new_n690_ = ~new_n688_ & ~new_n689_;
  assign new_n691_ = n11_ntk1 & ~new_n690_;
  assign new_n692_ = ~new_n232_ & ~new_n691_;
  assign new_n693_ = new_n224_ & new_n692_;
  assign new_n694_ = new_n686_ & ~new_n693_;
  assign new_n695_ = ~new_n686_ & new_n693_;
  assign new_n696_ = ~new_n694_ & ~new_n695_;
  assign new_n697_ = new_n246_ & new_n696_;
  assign new_n698_ = ~new_n687_ & ~new_n697_;
  assign new_n699_ = \o:~n68->n10  & new_n698_;
  assign new_n700_ = ~new_n228_ & ~new_n692_;
  assign new_n701_ = ~new_n223_ & ~new_n243_;
  assign new_n702_ = new_n700_ & new_n701_;
  assign new_n703_ = ~new_n700_ & ~new_n701_;
  assign new_n704_ = ~new_n702_ & ~new_n703_;
  assign new_n705_ = ~new_n228_ & ~new_n232_;
  assign new_n706_ = new_n691_ & new_n705_;
  assign new_n707_ = ~new_n691_ & ~new_n705_;
  assign new_n708_ = ~new_n706_ & ~new_n707_;
  assign new_n709_ = new_n704_ & new_n708_;
  assign new_n710_ = ~new_n215_ & ~new_n219_;
  assign new_n711_ = ~new_n223_ & ~new_n700_;
  assign new_n712_ = ~new_n243_ & ~new_n711_;
  assign new_n713_ = ~new_n710_ & ~new_n712_;
  assign new_n714_ = new_n710_ & new_n712_;
  assign new_n715_ = ~new_n713_ & ~new_n714_;
  assign new_n716_ = ~new_n236_ & ~new_n691_;
  assign new_n717_ = new_n715_ & new_n716_;
  assign new_n718_ = new_n709_ & new_n717_;
  assign new_n719_ = ~\i:n12_control_1  & ~n73_ntk1;
  assign new_n720_ = \i:n12_control_1  & ~n80_ntk1;
  assign new_n721_ = ~new_n719_ & ~new_n720_;
  assign new_n722_ = \i:n12_control_2  & ~new_n721_;
  assign new_n723_ = ~\i:n12_control_1  & ~n35_ntk1;
  assign new_n724_ = \i:n12_control_1  & ~n41_ntk1;
  assign new_n725_ = ~new_n723_ & ~new_n724_;
  assign new_n726_ = ~\i:n12_control_2  & ~new_n725_;
  assign new_n727_ = ~new_n722_ & ~new_n726_;
  assign new_n728_ = \i:n12_control_3  & ~new_n727_;
  assign new_n729_ = ~\i:n12_control_1  & ~n15_ntk1;
  assign new_n730_ = \i:n12_control_1  & ~n21_ntk1;
  assign new_n731_ = ~new_n729_ & ~new_n730_;
  assign new_n732_ = \i:n12_control_2  & ~new_n731_;
  assign new_n733_ = ~\i:n12_control_1  & ~n0_ntk1;
  assign new_n734_ = \i:n12_control_1  & ~n11_ntk1;
  assign new_n735_ = ~new_n733_ & ~new_n734_;
  assign new_n736_ = ~\i:n12_control_2  & ~new_n735_;
  assign new_n737_ = ~new_n732_ & ~new_n736_;
  assign new_n738_ = ~\i:n12_control_3  & ~new_n737_;
  assign new_n739_ = ~new_n728_ & ~new_n738_;
  assign new_n740_ = ~\i:n12_control_4  & ~new_n739_;
  assign new_n741_ = \i:n12_control_0  & new_n740_;
  assign new_n742_ = ~\i:n12_control_0  & ~new_n740_;
  assign new_n743_ = ~new_n741_ & ~new_n742_;
  assign new_n744_ = ~new_n677_ & ~new_n681_;
  assign new_n745_ = ~new_n642_ & new_n744_;
  assign new_n746_ = new_n644_ & ~new_n745_;
  assign new_n747_ = new_n743_ & ~new_n746_;
  assign new_n748_ = ~new_n506_ & ~new_n648_;
  assign new_n749_ = ~new_n747_ & ~new_n748_;
  assign new_n750_ = new_n747_ & new_n748_;
  assign new_n751_ = ~new_n749_ & ~new_n750_;
  assign new_n752_ = ~new_n677_ & new_n743_;
  assign new_n753_ = ~new_n638_ & ~new_n681_;
  assign new_n754_ = new_n752_ & ~new_n753_;
  assign new_n755_ = ~new_n752_ & new_n753_;
  assign new_n756_ = ~new_n754_ & ~new_n755_;
  assign new_n757_ = ~new_n751_ & new_n756_;
  assign new_n758_ = ~new_n648_ & new_n745_;
  assign new_n759_ = new_n650_ & ~new_n758_;
  assign new_n760_ = new_n743_ & ~new_n759_;
  assign new_n761_ = ~new_n374_ & ~new_n428_;
  assign new_n762_ = ~new_n760_ & ~new_n761_;
  assign new_n763_ = new_n760_ & new_n761_;
  assign new_n764_ = ~new_n762_ & ~new_n763_;
  assign new_n765_ = ~new_n638_ & ~new_n744_;
  assign new_n766_ = new_n743_ & ~new_n765_;
  assign new_n767_ = ~new_n584_ & ~new_n642_;
  assign new_n768_ = ~new_n766_ & ~new_n767_;
  assign new_n769_ = new_n766_ & new_n767_;
  assign new_n770_ = ~new_n768_ & ~new_n769_;
  assign new_n771_ = ~new_n764_ & ~new_n770_;
  assign new_n772_ = new_n757_ & new_n771_;
  assign new_n773_ = new_n718_ & ~new_n772_;
  assign new_n774_ = ~new_n718_ & new_n772_;
  assign new_n775_ = ~new_n773_ & ~new_n774_;
  assign new_n776_ = \o:~n56->n79  & new_n775_;
  assign new_n777_ = \o:n68->n10  & ~new_n698_;
  assign new_n778_ = ~new_n776_ & ~new_n777_;
  assign new_n779_ = ~new_n699_ & new_n778_;
  assign new_n780_ = \o:n56->n79  & ~new_n775_;
  assign new_n781_ = new_n716_ & ~new_n772_;
  assign new_n782_ = ~new_n716_ & new_n772_;
  assign new_n783_ = ~new_n781_ & ~new_n782_;
  assign new_n784_ = \o:~n56->n70  & new_n783_;
  assign new_n785_ = ~new_n693_ & ~new_n772_;
  assign new_n786_ = new_n693_ & new_n772_;
  assign new_n787_ = ~new_n785_ & ~new_n786_;
  assign new_n788_ = ~\o:~n56->n71  & new_n787_;
  assign new_n789_ = ~\o:n56->n71  & ~new_n787_;
  assign new_n790_ = ~new_n788_ & ~new_n789_;
  assign new_n791_ = ~new_n784_ & ~new_n790_;
  assign new_n792_ = ~new_n780_ & new_n791_;
  assign new_n793_ = ~new_n686_ & ~new_n718_;
  assign new_n794_ = new_n686_ & new_n718_;
  assign new_n795_ = ~new_n793_ & ~new_n794_;
  assign new_n796_ = \o:~n68->n79  & new_n795_;
  assign new_n797_ = \o:n68->n79  & ~new_n795_;
  assign new_n798_ = new_n246_ & ~new_n686_;
  assign new_n799_ = ~new_n687_ & ~new_n798_;
  assign new_n800_ = ~\o:~n68->n33  & ~new_n799_;
  assign new_n801_ = ~\o:n68->n33  & new_n799_;
  assign new_n802_ = ~new_n800_ & ~new_n801_;
  assign new_n803_ = ~new_n797_ & ~new_n802_;
  assign new_n804_ = ~new_n796_ & new_n803_;
  assign new_n805_ = ~new_n686_ & ~new_n704_;
  assign new_n806_ = new_n686_ & new_n704_;
  assign new_n807_ = ~new_n805_ & ~new_n806_;
  assign new_n808_ = ~\o:~n68->n39  & new_n807_;
  assign new_n809_ = ~\o:n68->n39  & ~new_n807_;
  assign new_n810_ = ~new_n808_ & ~new_n809_;
  assign new_n811_ = ~new_n686_ & ~new_n708_;
  assign new_n812_ = new_n686_ & new_n708_;
  assign new_n813_ = ~new_n811_ & ~new_n812_;
  assign new_n814_ = ~\o:~n68->n66  & new_n813_;
  assign new_n815_ = ~\o:n68->n66  & ~new_n813_;
  assign new_n816_ = ~new_n814_ & ~new_n815_;
  assign new_n817_ = ~new_n810_ & ~new_n816_;
  assign new_n818_ = new_n652_ & ~new_n704_;
  assign new_n819_ = ~new_n652_ & new_n704_;
  assign new_n820_ = ~new_n818_ & ~new_n819_;
  assign new_n821_ = ~\o:~n48->n39  & new_n820_;
  assign new_n822_ = ~\o:n48->n39  & ~new_n820_;
  assign new_n823_ = ~new_n821_ & ~new_n822_;
  assign new_n824_ = new_n652_ & ~new_n708_;
  assign new_n825_ = ~new_n652_ & new_n708_;
  assign new_n826_ = ~new_n824_ & ~new_n825_;
  assign new_n827_ = ~\o:~n48->n66  & new_n826_;
  assign new_n828_ = ~\o:n48->n66  & ~new_n826_;
  assign new_n829_ = ~new_n827_ & ~new_n828_;
  assign new_n830_ = ~new_n823_ & ~new_n829_;
  assign new_n831_ = ~new_n704_ & ~new_n770_;
  assign new_n832_ = new_n704_ & new_n770_;
  assign new_n833_ = ~new_n831_ & ~new_n832_;
  assign new_n834_ = \o:n42->n39  & ~new_n833_;
  assign new_n835_ = ~new_n716_ & ~new_n770_;
  assign new_n836_ = new_n716_ & new_n770_;
  assign new_n837_ = ~new_n835_ & ~new_n836_;
  assign new_n838_ = \o:~n42->n70  & new_n837_;
  assign new_n839_ = ~new_n684_ & ~new_n716_;
  assign new_n840_ = new_n684_ & new_n716_;
  assign new_n841_ = ~new_n839_ & ~new_n840_;
  assign new_n842_ = \o:~n77->n70  & new_n841_;
  assign new_n843_ = new_n684_ & ~new_n693_;
  assign new_n844_ = ~new_n684_ & new_n693_;
  assign new_n845_ = ~new_n843_ & ~new_n844_;
  assign new_n846_ = \o:n77->n71  & ~new_n845_;
  assign new_n847_ = ~new_n842_ & ~new_n846_;
  assign new_n848_ = \o:n77->n70  & ~new_n841_;
  assign new_n849_ = \o:~n77->n71  & new_n845_;
  assign new_n850_ = ~new_n848_ & ~new_n849_;
  assign new_n851_ = new_n847_ & new_n850_;
  assign new_n852_ = ~new_n838_ & new_n851_;
  assign new_n853_ = ~new_n834_ & new_n852_;
  assign new_n854_ = new_n693_ & ~new_n770_;
  assign new_n855_ = ~new_n693_ & new_n770_;
  assign new_n856_ = ~new_n854_ & ~new_n855_;
  assign new_n857_ = \o:n42->n71  & ~new_n856_;
  assign new_n858_ = \o:~n42->n39  & new_n833_;
  assign new_n859_ = ~new_n708_ & ~new_n770_;
  assign new_n860_ = new_n708_ & new_n770_;
  assign new_n861_ = ~new_n859_ & ~new_n860_;
  assign new_n862_ = \o:n42->n66  & ~new_n861_;
  assign new_n863_ = ~new_n858_ & ~new_n862_;
  assign new_n864_ = ~new_n857_ & new_n863_;
  assign new_n865_ = new_n853_ & new_n864_;
  assign new_n866_ = new_n830_ & new_n865_;
  assign new_n867_ = new_n817_ & new_n866_;
  assign new_n868_ = new_n804_ & new_n867_;
  assign new_n869_ = new_n792_ & new_n868_;
  assign new_n870_ = new_n779_ & new_n869_;
  assign new_n871_ = ~new_n718_ & ~new_n751_;
  assign new_n872_ = new_n718_ & new_n751_;
  assign new_n873_ = ~new_n871_ & ~new_n872_;
  assign new_n874_ = \o:~n9->n79  & new_n873_;
  assign new_n875_ = \o:n9->n79  & ~new_n873_;
  assign new_n876_ = ~new_n246_ & new_n652_;
  assign new_n877_ = new_n246_ & ~new_n652_;
  assign new_n878_ = ~new_n876_ & ~new_n877_;
  assign new_n879_ = ~\o:~n48->n33  & new_n878_;
  assign new_n880_ = ~\o:n48->n33  & ~new_n878_;
  assign new_n881_ = ~new_n879_ & ~new_n880_;
  assign new_n882_ = ~new_n875_ & ~new_n881_;
  assign new_n883_ = ~new_n874_ & new_n882_;
  assign new_n884_ = ~new_n246_ & new_n751_;
  assign new_n885_ = new_n246_ & ~new_n751_;
  assign new_n886_ = ~new_n884_ & ~new_n885_;
  assign new_n887_ = ~\o:~n9->n33  & ~new_n886_;
  assign new_n888_ = ~\o:n9->n33  & new_n886_;
  assign new_n889_ = ~new_n887_ & ~new_n888_;
  assign new_n890_ = ~new_n704_ & ~new_n751_;
  assign new_n891_ = new_n704_ & new_n751_;
  assign new_n892_ = ~new_n890_ & ~new_n891_;
  assign new_n893_ = ~\o:~n9->n39  & new_n892_;
  assign new_n894_ = ~\o:n9->n39  & ~new_n892_;
  assign new_n895_ = ~new_n893_ & ~new_n894_;
  assign new_n896_ = ~new_n889_ & ~new_n895_;
  assign new_n897_ = new_n883_ & new_n896_;
  assign new_n898_ = ~new_n716_ & ~new_n764_;
  assign new_n899_ = new_n716_ & new_n764_;
  assign new_n900_ = ~new_n898_ & ~new_n899_;
  assign new_n901_ = \o:n65->n70  & ~new_n900_;
  assign new_n902_ = \o:~n65->n70  & new_n900_;
  assign new_n903_ = ~new_n901_ & ~new_n902_;
  assign new_n904_ = ~new_n708_ & ~new_n764_;
  assign new_n905_ = new_n708_ & new_n764_;
  assign new_n906_ = ~new_n904_ & ~new_n905_;
  assign new_n907_ = \o:~n65->n66  & new_n906_;
  assign new_n908_ = \o:n65->n66  & ~new_n906_;
  assign new_n909_ = ~new_n907_ & ~new_n908_;
  assign new_n910_ = new_n903_ & new_n909_;
  assign new_n911_ = ~new_n718_ & ~new_n764_;
  assign new_n912_ = new_n718_ & new_n764_;
  assign new_n913_ = ~new_n911_ & ~new_n912_;
  assign new_n914_ = \o:~n65->n79  & new_n913_;
  assign new_n915_ = new_n693_ & ~new_n764_;
  assign new_n916_ = ~new_n693_ & new_n764_;
  assign new_n917_ = ~new_n915_ & ~new_n916_;
  assign new_n918_ = \o:~n65->n71  & new_n917_;
  assign new_n919_ = \o:n65->n79  & ~new_n913_;
  assign new_n920_ = ~new_n918_ & ~new_n919_;
  assign new_n921_ = ~new_n914_ & new_n920_;
  assign new_n922_ = \o:n65->n71  & ~new_n917_;
  assign new_n923_ = ~new_n246_ & new_n764_;
  assign new_n924_ = new_n246_ & ~new_n764_;
  assign new_n925_ = ~new_n923_ & ~new_n924_;
  assign new_n926_ = \o:~n65->n33  & ~new_n925_;
  assign new_n927_ = ~new_n922_ & ~new_n926_;
  assign new_n928_ = new_n921_ & new_n927_;
  assign new_n929_ = new_n910_ & new_n928_;
  assign new_n930_ = new_n897_ & new_n929_;
  assign new_n931_ = new_n708_ & ~new_n772_;
  assign new_n932_ = ~new_n708_ & new_n772_;
  assign new_n933_ = ~new_n931_ & ~new_n932_;
  assign new_n934_ = \o:n56->n66  & ~new_n933_;
  assign new_n935_ = \o:~n56->n66  & new_n933_;
  assign new_n936_ = ~new_n934_ & ~new_n935_;
  assign new_n937_ = new_n704_ & ~new_n772_;
  assign new_n938_ = ~new_n704_ & new_n772_;
  assign new_n939_ = ~new_n937_ & ~new_n938_;
  assign new_n940_ = \o:~n56->n39  & new_n939_;
  assign new_n941_ = \o:n56->n39  & ~new_n939_;
  assign new_n942_ = ~new_n940_ & ~new_n941_;
  assign new_n943_ = new_n936_ & new_n942_;
  assign new_n944_ = new_n715_ & ~new_n772_;
  assign new_n945_ = ~new_n715_ & new_n772_;
  assign new_n946_ = ~new_n944_ & ~new_n945_;
  assign new_n947_ = \o:n56->n4  & ~new_n946_;
  assign new_n948_ = ~new_n716_ & ~new_n751_;
  assign new_n949_ = new_n716_ & new_n751_;
  assign new_n950_ = ~new_n948_ & ~new_n949_;
  assign new_n951_ = \o:n9->n70  & ~new_n950_;
  assign new_n952_ = \o:~n9->n70  & new_n950_;
  assign new_n953_ = ~new_n951_ & ~new_n952_;
  assign new_n954_ = new_n693_ & ~new_n751_;
  assign new_n955_ = ~new_n693_ & new_n751_;
  assign new_n956_ = ~new_n954_ & ~new_n955_;
  assign new_n957_ = \o:n9->n71  & ~new_n956_;
  assign new_n958_ = \o:~n9->n71  & new_n956_;
  assign new_n959_ = ~new_n957_ & ~new_n958_;
  assign new_n960_ = new_n953_ & new_n959_;
  assign new_n961_ = new_n652_ & ~new_n716_;
  assign new_n962_ = ~new_n652_ & new_n716_;
  assign new_n963_ = ~new_n961_ & ~new_n962_;
  assign new_n964_ = ~\o:~n48->n70  & new_n963_;
  assign new_n965_ = ~\o:n48->n70  & ~new_n963_;
  assign new_n966_ = ~new_n964_ & ~new_n965_;
  assign new_n967_ = \o:~n42->n66  & new_n861_;
  assign new_n968_ = \o:n42->n70  & ~new_n837_;
  assign new_n969_ = ~new_n967_ & ~new_n968_;
  assign new_n970_ = ~new_n684_ & ~new_n708_;
  assign new_n971_ = new_n684_ & new_n708_;
  assign new_n972_ = ~new_n970_ & ~new_n971_;
  assign new_n973_ = \o:n77->n66  & ~new_n972_;
  assign new_n974_ = \o:~n77->n66  & new_n972_;
  assign new_n975_ = ~new_n973_ & ~new_n974_;
  assign new_n976_ = ~new_n684_ & ~new_n704_;
  assign new_n977_ = new_n684_ & new_n704_;
  assign new_n978_ = ~new_n976_ & ~new_n977_;
  assign new_n979_ = \o:n77->n39  & ~new_n978_;
  assign new_n980_ = \o:~n77->n39  & new_n978_;
  assign new_n981_ = ~\o:n65->n79  & ~\o:~n65->n79 ;
  assign new_n982_ = ~\o:~n65->n71  & new_n981_;
  assign new_n983_ = ~\o:~n65->n70  & ~\o:n65->n71 ;
  assign new_n984_ = ~\o:n65->n70  & new_n983_;
  assign new_n985_ = ~\o:~n65->n66  & new_n984_;
  assign new_n986_ = new_n982_ & new_n985_;
  assign new_n987_ = ~\o:n65->n66  & new_n986_;
  assign new_n988_ = ~\o:~n65->n39  & new_n987_;
  assign new_n989_ = ~\o:n65->n39  & new_n988_;
  assign new_n990_ = \o:~n65->n33  & ~new_n989_;
  assign new_n991_ = ~\o:n68->n4  & ~\o:~n68->n4 ;
  assign new_n992_ = ~\o:n65->n4  & ~\o:~n65->n4 ;
  assign new_n993_ = new_n991_ & new_n992_;
  assign new_n994_ = ~\o:~n9->n4  & new_n993_;
  assign new_n995_ = ~\o:n56->n4  & ~\o:~n56->n4 ;
  assign new_n996_ = ~\o:~n48->n4  & new_n995_;
  assign new_n997_ = ~\o:n48->n4  & new_n996_;
  assign new_n998_ = new_n994_ & new_n997_;
  assign new_n999_ = \o:n9->n4  & ~new_n998_;
  assign new_n1000_ = ~\o:n48->n10  & ~\o:~n48->n10 ;
  assign new_n1001_ = ~\o:n68->n10  & ~\o:~n68->n10 ;
  assign new_n1002_ = ~\o:n65->n10  & ~\o:~n65->n10 ;
  assign new_n1003_ = ~\o:n56->n10  & ~\o:~n56->n10 ;
  assign new_n1004_ = new_n1002_ & new_n1003_;
  assign new_n1005_ = \o:~n48->n10  & ~new_n1004_;
  assign new_n1006_ = new_n1001_ & ~new_n1005_;
  assign new_n1007_ = ~new_n1000_ & ~new_n1006_;
  assign new_n1008_ = ~new_n999_ & ~new_n1007_;
  assign new_n1009_ = new_n1001_ & new_n1002_;
  assign new_n1010_ = ~\o:~n9->n10  & new_n1009_;
  assign new_n1011_ = ~\o:~n48->n10  & new_n1003_;
  assign new_n1012_ = ~\o:n48->n10  & new_n1011_;
  assign new_n1013_ = new_n1010_ & new_n1012_;
  assign new_n1014_ = \o:n9->n10  & ~new_n1013_;
  assign new_n1015_ = new_n1008_ & ~new_n1014_;
  assign new_n1016_ = ~new_n990_ & new_n1015_;
  assign new_n1017_ = ~\o:~n56->n70  & ~\o:n65->n70 ;
  assign new_n1018_ = ~\o:n77->n70  & ~\o:~n77->n70 ;
  assign new_n1019_ = ~\o:~n68->n70  & new_n1018_;
  assign new_n1020_ = ~\o:~n65->n70  & ~\o:n68->n70 ;
  assign new_n1021_ = new_n1019_ & new_n1020_;
  assign new_n1022_ = new_n1017_ & new_n1021_;
  assign new_n1023_ = ~\o:n56->n70  & new_n1022_;
  assign new_n1024_ = ~\o:~n48->n70  & new_n1023_;
  assign new_n1025_ = ~\o:n48->n70  & new_n1024_;
  assign new_n1026_ = \o:~n42->n70  & ~new_n1025_;
  assign new_n1027_ = ~\o:n56->n79  & ~\o:~n56->n79 ;
  assign new_n1028_ = ~\o:~n56->n71  & new_n1027_;
  assign new_n1029_ = ~\o:~n56->n66  & ~\o:n56->n70 ;
  assign new_n1030_ = ~\o:~n56->n70  & ~\o:n56->n71 ;
  assign new_n1031_ = new_n1029_ & new_n1030_;
  assign new_n1032_ = new_n1028_ & new_n1031_;
  assign new_n1033_ = ~\o:n56->n66  & new_n1032_;
  assign new_n1034_ = ~\o:~n56->n39  & new_n1033_;
  assign new_n1035_ = ~\o:n56->n39  & new_n1034_;
  assign new_n1036_ = \o:~n56->n33  & ~new_n1035_;
  assign new_n1037_ = ~\o:n68->n79  & ~\o:~n68->n79 ;
  assign new_n1038_ = ~\o:~n68->n71  & new_n1037_;
  assign new_n1039_ = ~\o:~n68->n70  & ~\o:n68->n71 ;
  assign new_n1040_ = ~\o:n68->n70  & new_n1039_;
  assign new_n1041_ = ~\o:~n68->n66  & new_n1040_;
  assign new_n1042_ = new_n1038_ & new_n1041_;
  assign new_n1043_ = ~\o:n68->n66  & new_n1042_;
  assign new_n1044_ = ~\o:~n68->n39  & new_n1043_;
  assign new_n1045_ = \o:n68->n39  & ~new_n1044_;
  assign new_n1046_ = \o:n68->n66  & ~new_n1042_;
  assign new_n1047_ = ~new_n1045_ & ~new_n1046_;
  assign new_n1048_ = ~new_n1036_ & new_n1047_;
  assign new_n1049_ = ~new_n1026_ & new_n1048_;
  assign new_n1050_ = new_n1016_ & new_n1049_;
  assign new_n1051_ = ~\o:n56->n33  & ~\o:~n56->n33 ;
  assign new_n1052_ = new_n1035_ & new_n1051_;
  assign new_n1053_ = \o:~n56->n10  & ~new_n1052_;
  assign new_n1054_ = ~\o:n56->n10  & ~new_n1053_;
  assign new_n1055_ = ~\o:n56->n39  & ~\o:~n56->n39 ;
  assign new_n1056_ = new_n1051_ & new_n1055_;
  assign new_n1057_ = ~\o:n56->n70  & ~\o:~n56->n70 ;
  assign new_n1058_ = ~\o:n56->n66  & ~\o:~n56->n66 ;
  assign new_n1059_ = new_n1057_ & new_n1058_;
  assign new_n1060_ = ~\o:n56->n71  & new_n1028_;
  assign new_n1061_ = new_n1059_ & new_n1060_;
  assign new_n1062_ = ~\o:~n56->n10  & new_n1061_;
  assign new_n1063_ = new_n1056_ & new_n1062_;
  assign new_n1064_ = ~new_n1054_ & ~new_n1063_;
  assign new_n1065_ = new_n1050_ & ~new_n1064_;
  assign new_n1066_ = ~\o:n68->n66  & new_n1041_;
  assign new_n1067_ = ~\o:~n68->n71  & new_n1066_;
  assign new_n1068_ = \o:~n68->n39  & ~new_n1067_;
  assign new_n1069_ = ~\o:n9->n39  & ~\o:n42->n39 ;
  assign new_n1070_ = ~\o:n48->n39  & ~\o:~n48->n39 ;
  assign new_n1071_ = ~\o:n68->n39  & ~\o:~n68->n39 ;
  assign new_n1072_ = new_n1070_ & new_n1071_;
  assign new_n1073_ = new_n1069_ & new_n1072_;
  assign new_n1074_ = ~\o:n65->n39  & new_n1055_;
  assign new_n1075_ = ~\o:n77->n39  & ~\o:~n77->n39 ;
  assign new_n1076_ = new_n1074_ & new_n1075_;
  assign new_n1077_ = ~\o:~n65->n39  & new_n1076_;
  assign new_n1078_ = new_n1073_ & new_n1077_;
  assign new_n1079_ = \o:~n9->n39  & ~new_n1078_;
  assign new_n1080_ = ~new_n1068_ & ~new_n1079_;
  assign new_n1081_ = ~\o:n65->n70  & ~\o:~n65->n70 ;
  assign new_n1082_ = ~\o:n65->n71  & new_n982_;
  assign new_n1083_ = new_n1081_ & new_n1082_;
  assign new_n1084_ = \o:~n65->n66  & ~new_n1083_;
  assign new_n1085_ = \o:~n56->n4  & ~new_n1061_;
  assign new_n1086_ = new_n1028_ & new_n1030_;
  assign new_n1087_ = ~new_n1029_ & ~new_n1086_;
  assign new_n1088_ = ~\o:n65->n39  & ~\o:~n65->n39 ;
  assign new_n1089_ = ~\o:n65->n66  & ~\o:~n65->n66 ;
  assign new_n1090_ = ~\o:n65->n70  & new_n1089_;
  assign new_n1091_ = new_n1088_ & new_n1090_;
  assign new_n1092_ = \o:n65->n33  & ~new_n1091_;
  assign new_n1093_ = ~new_n1087_ & ~new_n1092_;
  assign new_n1094_ = ~new_n1085_ & new_n1093_;
  assign new_n1095_ = ~new_n1084_ & new_n1094_;
  assign new_n1096_ = new_n1080_ & new_n1095_;
  assign new_n1097_ = ~\o:n77->n71  & ~\o:~n77->n71 ;
  assign new_n1098_ = ~\o:n56->n71  & ~\o:~n56->n71 ;
  assign new_n1099_ = ~\o:n65->n71  & new_n1098_;
  assign new_n1100_ = new_n1097_ & new_n1099_;
  assign new_n1101_ = ~\o:~n65->n71  & ~\o:n68->n71 ;
  assign new_n1102_ = new_n1100_ & new_n1101_;
  assign new_n1103_ = \o:~n9->n71  & ~new_n1102_;
  assign new_n1104_ = ~\o:~n48->n79  & new_n1027_;
  assign new_n1105_ = new_n981_ & new_n1104_;
  assign new_n1106_ = \o:n48->n79  & ~new_n1105_;
  assign new_n1107_ = new_n981_ & new_n1027_;
  assign new_n1108_ = \o:~n48->n79  & ~new_n1107_;
  assign new_n1109_ = ~\o:~n9->n79  & ~new_n1108_;
  assign new_n1110_ = ~new_n1106_ & new_n1109_;
  assign new_n1111_ = new_n981_ & new_n1037_;
  assign new_n1112_ = ~\o:n48->n79  & new_n1104_;
  assign new_n1113_ = new_n1111_ & new_n1112_;
  assign new_n1114_ = ~new_n1110_ & ~new_n1113_;
  assign new_n1115_ = ~new_n1103_ & ~new_n1114_;
  assign new_n1116_ = new_n1058_ & new_n1089_;
  assign new_n1117_ = ~\o:n48->n66  & ~\o:~n48->n66 ;
  assign new_n1118_ = ~\o:n42->n66  & ~\o:~n42->n66 ;
  assign new_n1119_ = new_n1117_ & new_n1118_;
  assign new_n1120_ = new_n1116_ & new_n1119_;
  assign new_n1121_ = \o:~n6->n66  & ~new_n1120_;
  assign new_n1122_ = ~\o:n56->n39  & new_n1070_;
  assign new_n1123_ = ~\o:~n65->n39  & new_n1071_;
  assign new_n1124_ = ~\o:n65->n39  & new_n1123_;
  assign new_n1125_ = ~\o:~n56->n39  & new_n1124_;
  assign new_n1126_ = ~new_n1122_ & ~new_n1125_;
  assign new_n1127_ = ~new_n1121_ & ~new_n1126_;
  assign new_n1128_ = ~\o:n6->n66  & ~\o:~n6->n66 ;
  assign new_n1129_ = ~\o:n9->n66  & ~\o:~n9->n66 ;
  assign new_n1130_ = ~\o:n68->n66  & ~\o:~n68->n66 ;
  assign new_n1131_ = ~\o:n77->n66  & ~\o:~n77->n66 ;
  assign new_n1132_ = new_n1130_ & new_n1131_;
  assign new_n1133_ = new_n1129_ & new_n1132_;
  assign new_n1134_ = ~new_n1128_ & ~new_n1133_;
  assign new_n1135_ = ~\o:~n68->n66  & new_n1131_;
  assign new_n1136_ = ~\o:~n65->n66  & ~\o:n68->n66 ;
  assign new_n1137_ = new_n1135_ & new_n1136_;
  assign new_n1138_ = ~\o:n65->n66  & new_n1137_;
  assign new_n1139_ = \o:~n56->n66  & ~new_n1138_;
  assign new_n1140_ = ~new_n1134_ & ~new_n1139_;
  assign new_n1141_ = new_n1127_ & new_n1140_;
  assign new_n1142_ = new_n1115_ & new_n1141_;
  assign new_n1143_ = ~\o:~n48->n33  & new_n1051_;
  assign new_n1144_ = ~\o:n65->n33  & ~\o:~n65->n33 ;
  assign new_n1145_ = new_n1143_ & new_n1144_;
  assign new_n1146_ = \o:n48->n33  & ~new_n1145_;
  assign new_n1147_ = new_n1051_ & new_n1144_;
  assign new_n1148_ = \o:~n48->n33  & ~new_n1147_;
  assign new_n1149_ = ~\o:~n9->n33  & ~new_n1148_;
  assign new_n1150_ = ~new_n1146_ & new_n1149_;
  assign new_n1151_ = ~\o:n68->n33  & ~\o:~n68->n33 ;
  assign new_n1152_ = new_n1144_ & new_n1151_;
  assign new_n1153_ = ~\o:n48->n33  & new_n1143_;
  assign new_n1154_ = new_n1152_ & new_n1153_;
  assign new_n1155_ = ~new_n1150_ & ~new_n1154_;
  assign new_n1156_ = \o:~n56->n70  & \o:n65->n70 ;
  assign new_n1157_ = ~new_n1017_ & ~new_n1021_;
  assign new_n1158_ = ~new_n1156_ & ~new_n1157_;
  assign new_n1159_ = ~\o:~n9->n71  & ~\o:~n42->n71 ;
  assign new_n1160_ = ~\o:n48->n71  & ~\o:~n48->n71 ;
  assign new_n1161_ = ~\o:n9->n71  & ~\o:n42->n71 ;
  assign new_n1162_ = ~\o:~n68->n71  & new_n1161_;
  assign new_n1163_ = new_n1160_ & new_n1162_;
  assign new_n1164_ = ~new_n1159_ & ~new_n1163_;
  assign new_n1165_ = new_n1158_ & ~new_n1164_;
  assign new_n1166_ = ~new_n1155_ & new_n1165_;
  assign new_n1167_ = new_n1142_ & new_n1166_;
  assign new_n1168_ = new_n1096_ & new_n1167_;
  assign new_n1169_ = ~\o:n56->n70  & new_n1055_;
  assign new_n1170_ = new_n1058_ & new_n1086_;
  assign new_n1171_ = new_n1169_ & new_n1170_;
  assign new_n1172_ = \o:n56->n33  & ~new_n1171_;
  assign new_n1173_ = ~\o:n65->n66  & new_n985_;
  assign new_n1174_ = ~\o:~n65->n71  & new_n1173_;
  assign new_n1175_ = \o:~n65->n39  & ~new_n1174_;
  assign new_n1176_ = ~new_n1172_ & ~new_n1175_;
  assign new_n1177_ = new_n1038_ & new_n1039_;
  assign new_n1178_ = \o:n68->n70  & ~new_n1177_;
  assign new_n1179_ = ~\o:n68->n71  & new_n1038_;
  assign new_n1180_ = \o:~n68->n70  & ~new_n1179_;
  assign new_n1181_ = ~new_n1178_ & ~new_n1180_;
  assign new_n1182_ = new_n1018_ & new_n1097_;
  assign new_n1183_ = new_n1131_ & new_n1182_;
  assign new_n1184_ = \o:~n77->n39  & ~new_n1183_;
  assign new_n1185_ = new_n1181_ & ~new_n1184_;
  assign new_n1186_ = new_n993_ & new_n997_;
  assign new_n1187_ = \o:~n9->n4  & ~new_n1186_;
  assign new_n1188_ = new_n1009_ & new_n1012_;
  assign new_n1189_ = \o:~n9->n10  & ~new_n1188_;
  assign new_n1190_ = ~new_n1187_ & ~new_n1189_;
  assign new_n1191_ = new_n1185_ & new_n1190_;
  assign new_n1192_ = \o:~n56->n66  & \o:n56->n70 ;
  assign new_n1193_ = new_n982_ & new_n983_;
  assign new_n1194_ = \o:n65->n70  & ~new_n1193_;
  assign new_n1195_ = \o:~n65->n70  & ~new_n1082_;
  assign new_n1196_ = ~new_n1194_ & ~new_n1195_;
  assign new_n1197_ = new_n1071_ & new_n1151_;
  assign new_n1198_ = new_n1001_ & new_n1197_;
  assign new_n1199_ = ~new_n991_ & ~new_n1198_;
  assign new_n1200_ = new_n1196_ & ~new_n1199_;
  assign new_n1201_ = ~new_n1192_ & new_n1200_;
  assign new_n1202_ = new_n1191_ & new_n1201_;
  assign new_n1203_ = new_n1176_ & new_n1202_;
  assign new_n1204_ = ~\o:n68->n71  & ~\o:~n68->n71 ;
  assign new_n1205_ = ~\o:~n65->n71  & new_n1204_;
  assign new_n1206_ = ~\o:n65->n71  & new_n1205_;
  assign new_n1207_ = \o:~n56->n71  & ~new_n1206_;
  assign new_n1208_ = ~\o:~n56->n71  & new_n1206_;
  assign new_n1209_ = new_n1097_ & new_n1208_;
  assign new_n1210_ = ~new_n1160_ & ~new_n1209_;
  assign new_n1211_ = ~new_n1207_ & ~new_n1210_;
  assign new_n1212_ = new_n1055_ & new_n1123_;
  assign new_n1213_ = ~new_n1075_ & ~new_n1212_;
  assign new_n1214_ = \o:~n56->n39  & ~new_n1124_;
  assign new_n1215_ = ~\o:n56->n39  & new_n1075_;
  assign new_n1216_ = ~new_n1070_ & ~new_n1215_;
  assign new_n1217_ = ~new_n1214_ & ~new_n1216_;
  assign new_n1218_ = ~new_n1213_ & new_n1217_;
  assign new_n1219_ = ~\o:n65->n70  & new_n1057_;
  assign new_n1220_ = ~\o:n42->n70  & ~\o:~n48->n70 ;
  assign new_n1221_ = ~new_n1219_ & ~new_n1220_;
  assign new_n1222_ = new_n1218_ & ~new_n1221_;
  assign new_n1223_ = new_n1211_ & new_n1222_;
  assign new_n1224_ = new_n1203_ & new_n1223_;
  assign new_n1225_ = new_n1168_ & new_n1224_;
  assign new_n1226_ = ~\o:n48->n79  & ~\o:~n48->n79 ;
  assign new_n1227_ = ~\o:~n48->n71  & new_n1226_;
  assign new_n1228_ = ~\o:n48->n71  & new_n1227_;
  assign new_n1229_ = \o:n48->n79  & \o:~n48->n79 ;
  assign new_n1230_ = ~\o:~n48->n70  & ~new_n1229_;
  assign new_n1231_ = ~new_n1228_ & ~new_n1230_;
  assign new_n1232_ = ~\o:~n48->n70  & ~\o:n48->n71 ;
  assign new_n1233_ = new_n1227_ & new_n1232_;
  assign new_n1234_ = \o:n48->n70  & ~new_n1233_;
  assign new_n1235_ = new_n1003_ & new_n1056_;
  assign new_n1236_ = ~new_n995_ & ~new_n1235_;
  assign new_n1237_ = ~new_n1234_ & ~new_n1236_;
  assign new_n1238_ = ~new_n1231_ & new_n1237_;
  assign new_n1239_ = ~\o:n42->n70  & ~\o:~n42->n70 ;
  assign new_n1240_ = ~\o:n42->n71  & ~\o:~n42->n71 ;
  assign new_n1241_ = new_n1239_ & new_n1240_;
  assign new_n1242_ = new_n1118_ & new_n1241_;
  assign new_n1243_ = ~\o:~n42->n39  & new_n1242_;
  assign new_n1244_ = ~\o:n42->n39  & new_n1243_;
  assign new_n1245_ = new_n1117_ & new_n1233_;
  assign new_n1246_ = ~\o:~n48->n33  & new_n1070_;
  assign new_n1247_ = ~\o:n48->n70  & new_n1246_;
  assign new_n1248_ = new_n1245_ & new_n1247_;
  assign new_n1249_ = \o:n48->n33  & ~new_n1248_;
  assign new_n1250_ = ~new_n1244_ & ~new_n1249_;
  assign new_n1251_ = ~\o:n6->n71  & ~\o:~n6->n71 ;
  assign new_n1252_ = \o:n42->n70  & \o:~n42->n70 ;
  assign new_n1253_ = \o:n48->n71  & \o:~n48->n71 ;
  assign new_n1254_ = ~new_n1252_ & ~new_n1253_;
  assign new_n1255_ = \o:n65->n33  & \o:~n65->n33 ;
  assign new_n1256_ = \o:n65->n71  & \o:~n65->n71 ;
  assign new_n1257_ = ~new_n1255_ & ~new_n1256_;
  assign new_n1258_ = \o:n68->n33  & \o:~n68->n33 ;
  assign new_n1259_ = \o:n56->n79  & \o:~n56->n79 ;
  assign new_n1260_ = ~new_n1258_ & ~new_n1259_;
  assign new_n1261_ = new_n1257_ & new_n1260_;
  assign new_n1262_ = new_n1254_ & new_n1261_;
  assign new_n1263_ = new_n1251_ & new_n1262_;
  assign new_n1264_ = \o:n42->n66  & \o:~n42->n66 ;
  assign new_n1265_ = ~\o:n6->n4  & ~new_n1264_;
  assign new_n1266_ = ~\o:~n6->n4  & new_n1265_;
  assign new_n1267_ = \o:n9->n79  & \o:~n9->n79 ;
  assign new_n1268_ = ~\o:n6->n33  & ~\o:~n6->n33 ;
  assign new_n1269_ = ~\o:n6->n39  & ~\o:~n6->n39 ;
  assign new_n1270_ = ~\o:~n6->n10  & new_n1269_;
  assign new_n1271_ = new_n1268_ & new_n1270_;
  assign new_n1272_ = ~new_n1267_ & new_n1271_;
  assign new_n1273_ = new_n1266_ & new_n1272_;
  assign new_n1274_ = new_n1263_ & new_n1273_;
  assign new_n1275_ = new_n1250_ & new_n1274_;
  assign new_n1276_ = new_n1238_ & new_n1275_;
  assign new_n1277_ = ~\o:n9->n79  & ~\o:~n9->n79 ;
  assign new_n1278_ = ~\o:~n9->n71  & new_n1277_;
  assign new_n1279_ = \o:~n9->n70  & ~new_n1278_;
  assign new_n1280_ = ~\o:n9->n71  & new_n1277_;
  assign new_n1281_ = ~\o:~n9->n70  & new_n1277_;
  assign new_n1282_ = \o:n9->n71  & ~new_n1281_;
  assign new_n1283_ = ~\o:~n9->n71  & ~new_n1282_;
  assign new_n1284_ = ~new_n1280_ & ~new_n1283_;
  assign new_n1285_ = ~\o:n42->n71  & new_n1239_;
  assign new_n1286_ = \o:~n42->n66  & ~new_n1285_;
  assign new_n1287_ = new_n1075_ & new_n1183_;
  assign new_n1288_ = ~new_n1286_ & ~new_n1287_;
  assign new_n1289_ = ~new_n1284_ & new_n1288_;
  assign new_n1290_ = ~new_n1279_ & new_n1289_;
  assign new_n1291_ = ~\o:n56->n71  & new_n1027_;
  assign new_n1292_ = \o:~n56->n71  & ~new_n1291_;
  assign new_n1293_ = \o:n68->n39  & \o:~n68->n39 ;
  assign new_n1294_ = \o:n68->n10  & \o:~n68->n10 ;
  assign new_n1295_ = \o:n9->n39  & \o:n42->n39 ;
  assign new_n1296_ = ~new_n1294_ & ~new_n1295_;
  assign new_n1297_ = \o:~n42->n71  & \o:~n77->n71 ;
  assign new_n1298_ = \o:~n42->n39  & \o:~n77->n39 ;
  assign new_n1299_ = ~new_n1297_ & ~new_n1298_;
  assign new_n1300_ = new_n1296_ & new_n1299_;
  assign new_n1301_ = ~new_n1293_ & new_n1300_;
  assign new_n1302_ = \o:n65->n4  & \o:~n65->n4 ;
  assign new_n1303_ = \o:n68->n71  & \o:~n68->n71 ;
  assign new_n1304_ = \o:n68->n79  & \o:~n68->n79 ;
  assign new_n1305_ = ~new_n1303_ & ~new_n1304_;
  assign new_n1306_ = ~new_n1302_ & new_n1305_;
  assign new_n1307_ = new_n1301_ & new_n1306_;
  assign new_n1308_ = \o:n65->n10  & \o:~n65->n10 ;
  assign new_n1309_ = \o:n77->n71  & \o:~n77->n71 ;
  assign new_n1310_ = \o:n77->n70  & \o:~n77->n70 ;
  assign new_n1311_ = ~new_n1309_ & ~new_n1310_;
  assign new_n1312_ = ~new_n1308_ & new_n1311_;
  assign new_n1313_ = ~\o:n6->n79  & ~\o:~n6->n79 ;
  assign new_n1314_ = ~\o:n6->n10  & new_n1313_;
  assign new_n1315_ = \o:n65->n79  & \o:~n65->n79 ;
  assign new_n1316_ = \o:n56->n33  & \o:~n56->n33 ;
  assign new_n1317_ = ~new_n1315_ & ~new_n1316_;
  assign new_n1318_ = new_n1314_ & new_n1317_;
  assign new_n1319_ = new_n1312_ & new_n1318_;
  assign new_n1320_ = \o:n68->n4  & \o:~n68->n4 ;
  assign new_n1321_ = \o:n77->n66  & \o:~n77->n66 ;
  assign new_n1322_ = ~new_n1320_ & ~new_n1321_;
  assign new_n1323_ = \o:n9->n71  & \o:n42->n71 ;
  assign new_n1324_ = \o:n48->n39  & \o:~n48->n39 ;
  assign new_n1325_ = ~new_n1323_ & ~new_n1324_;
  assign new_n1326_ = new_n1322_ & new_n1325_;
  assign new_n1327_ = \o:n42->n66  & ~new_n1241_;
  assign new_n1328_ = ~\o:n6->n70  & ~\o:~n6->n70 ;
  assign new_n1329_ = \o:n6->n66  & \o:~n6->n66 ;
  assign new_n1330_ = new_n1328_ & ~new_n1329_;
  assign new_n1331_ = \o:n6->n70  & \o:~n6->n70 ;
  assign new_n1332_ = new_n1128_ & ~new_n1331_;
  assign new_n1333_ = ~new_n1330_ & ~new_n1332_;
  assign new_n1334_ = ~new_n1327_ & ~new_n1333_;
  assign new_n1335_ = new_n1326_ & new_n1334_;
  assign new_n1336_ = new_n1319_ & new_n1335_;
  assign new_n1337_ = new_n1307_ & new_n1336_;
  assign new_n1338_ = ~new_n1292_ & new_n1337_;
  assign new_n1339_ = new_n1290_ & new_n1338_;
  assign new_n1340_ = new_n1276_ & new_n1339_;
  assign new_n1341_ = new_n1225_ & new_n1340_;
  assign new_n1342_ = \o:n68->n33  & ~new_n1177_;
  assign new_n1343_ = ~\o:n68->n70  & ~\o:~n68->n70 ;
  assign new_n1344_ = new_n1179_ & new_n1343_;
  assign new_n1345_ = new_n1130_ & new_n1344_;
  assign new_n1346_ = \o:~n68->n4  & ~new_n1345_;
  assign new_n1347_ = new_n992_ & new_n996_;
  assign new_n1348_ = \o:n48->n4  & ~new_n1347_;
  assign new_n1349_ = new_n1002_ & new_n1011_;
  assign new_n1350_ = \o:n48->n10  & ~new_n1349_;
  assign new_n1351_ = ~new_n1018_ & ~new_n1097_;
  assign new_n1352_ = ~\o:~n77->n66  & ~new_n1351_;
  assign new_n1353_ = ~new_n1182_ & ~new_n1352_;
  assign new_n1354_ = ~new_n1350_ & ~new_n1353_;
  assign new_n1355_ = ~new_n1348_ & new_n1354_;
  assign new_n1356_ = ~new_n1346_ & new_n1355_;
  assign new_n1357_ = ~new_n1342_ & new_n1356_;
  assign new_n1358_ = \o:n65->n33  & ~new_n1193_;
  assign new_n1359_ = ~\o:~n77->n39  & new_n1183_;
  assign new_n1360_ = \o:n77->n39  & ~new_n1359_;
  assign new_n1361_ = \o:~n68->n66  & ~new_n1344_;
  assign new_n1362_ = new_n1055_ & new_n1088_;
  assign new_n1363_ = ~\o:~n9->n39  & ~\o:n77->n39 ;
  assign new_n1364_ = new_n1362_ & new_n1363_;
  assign new_n1365_ = new_n1073_ & new_n1364_;
  assign new_n1366_ = \o:~n42->n39  & ~new_n1365_;
  assign new_n1367_ = ~new_n1361_ & ~new_n1366_;
  assign new_n1368_ = ~new_n1360_ & new_n1367_;
  assign new_n1369_ = ~new_n1358_ & new_n1368_;
  assign new_n1370_ = new_n1357_ & new_n1369_;
  assign new_n1371_ = new_n1129_ & new_n1280_;
  assign new_n1372_ = ~\o:~n9->n71  & new_n1371_;
  assign new_n1373_ = ~\o:n9->n70  & ~\o:~n9->n70 ;
  assign new_n1374_ = ~\o:n9->n33  & ~\o:~n9->n33 ;
  assign new_n1375_ = ~\o:n9->n39  & ~\o:~n9->n39 ;
  assign new_n1376_ = new_n1374_ & new_n1375_;
  assign new_n1377_ = new_n1373_ & new_n1376_;
  assign new_n1378_ = new_n1372_ & new_n1377_;
  assign new_n1379_ = ~\o:n9->n10  & new_n1378_;
  assign new_n1380_ = ~\o:~n9->n10  & new_n1379_;
  assign new_n1381_ = ~\o:~n9->n4  & new_n1380_;
  assign new_n1382_ = ~\o:n9->n4  & new_n1381_;
  assign new_n1383_ = ~\o:n68->n70  & new_n1130_;
  assign new_n1384_ = new_n1071_ & new_n1383_;
  assign new_n1385_ = \o:n68->n33  & ~new_n1384_;
  assign new_n1386_ = new_n1083_ & new_n1089_;
  assign new_n1387_ = \o:~n65->n4  & ~new_n1386_;
  assign new_n1388_ = new_n1088_ & new_n1144_;
  assign new_n1389_ = new_n1002_ & new_n1388_;
  assign new_n1390_ = ~new_n992_ & ~new_n1389_;
  assign new_n1391_ = ~\o:n56->n66  & new_n1031_;
  assign new_n1392_ = ~\o:~n56->n71  & new_n1391_;
  assign new_n1393_ = \o:~n56->n39  & ~new_n1392_;
  assign new_n1394_ = ~new_n1390_ & ~new_n1393_;
  assign new_n1395_ = ~new_n1387_ & new_n1394_;
  assign new_n1396_ = ~new_n1385_ & new_n1395_;
  assign new_n1397_ = ~\o:n65->n71  & ~\o:~n65->n71 ;
  assign new_n1398_ = new_n1098_ & new_n1397_;
  assign new_n1399_ = ~\o:~n9->n71  & ~\o:n68->n71 ;
  assign new_n1400_ = ~\o:n77->n71  & new_n1399_;
  assign new_n1401_ = new_n1398_ & new_n1400_;
  assign new_n1402_ = \o:~n42->n71  & ~new_n1401_;
  assign new_n1403_ = new_n1160_ & new_n1208_;
  assign new_n1404_ = \o:n56->n71  & ~new_n1403_;
  assign new_n1405_ = ~new_n1402_ & ~new_n1404_;
  assign new_n1406_ = ~\o:n65->n66  & new_n1058_;
  assign new_n1407_ = new_n1117_ & new_n1406_;
  assign new_n1408_ = new_n1137_ & new_n1407_;
  assign new_n1409_ = \o:n42->n66  & ~new_n1408_;
  assign new_n1410_ = ~\o:n48->n70  & ~\o:~n48->n70 ;
  assign new_n1411_ = new_n1021_ & new_n1410_;
  assign new_n1412_ = \o:n42->n70  & ~new_n1411_;
  assign new_n1413_ = ~new_n1409_ & ~new_n1412_;
  assign new_n1414_ = \o:n65->n66  & ~new_n1137_;
  assign new_n1415_ = ~\o:n68->n70  & new_n1019_;
  assign new_n1416_ = new_n1373_ & new_n1415_;
  assign new_n1417_ = ~new_n1328_ & ~new_n1416_;
  assign new_n1418_ = ~new_n1414_ & ~new_n1417_;
  assign new_n1419_ = new_n1057_ & new_n1081_;
  assign new_n1420_ = new_n1239_ & new_n1410_;
  assign new_n1421_ = new_n1419_ & new_n1420_;
  assign new_n1422_ = \o:~n6->n70  & ~new_n1421_;
  assign new_n1423_ = ~\o:~n68->n70  & new_n1020_;
  assign new_n1424_ = \o:~n48->n70  & ~new_n1423_;
  assign new_n1425_ = ~new_n1422_ & ~new_n1424_;
  assign new_n1426_ = ~\o:~n68->n66  & new_n1136_;
  assign new_n1427_ = new_n1406_ & new_n1426_;
  assign new_n1428_ = \o:~n48->n66  & ~new_n1427_;
  assign new_n1429_ = new_n1425_ & ~new_n1428_;
  assign new_n1430_ = new_n1418_ & new_n1429_;
  assign new_n1431_ = new_n1413_ & new_n1430_;
  assign new_n1432_ = new_n1405_ & new_n1431_;
  assign new_n1433_ = new_n1396_ & new_n1432_;
  assign new_n1434_ = ~new_n1382_ & new_n1433_;
  assign new_n1435_ = new_n1370_ & new_n1434_;
  assign new_n1436_ = new_n1341_ & new_n1435_;
  assign new_n1437_ = new_n1065_ & new_n1436_;
  assign new_n1438_ = new_n1415_ & new_n1421_;
  assign new_n1439_ = \o:n9->n70  & ~new_n1438_;
  assign new_n1440_ = \o:n48->n4  & \o:~n48->n4 ;
  assign new_n1441_ = ~\o:n48->n33  & ~\o:~n48->n33 ;
  assign new_n1442_ = new_n1070_ & new_n1441_;
  assign new_n1443_ = new_n1228_ & new_n1410_;
  assign new_n1444_ = new_n1117_ & new_n1443_;
  assign new_n1445_ = new_n1442_ & new_n1444_;
  assign new_n1446_ = ~\o:~n48->n10  & new_n1445_;
  assign new_n1447_ = \o:n48->n10  & ~new_n1446_;
  assign new_n1448_ = ~new_n1440_ & ~new_n1447_;
  assign new_n1449_ = ~new_n1439_ & new_n1448_;
  assign new_n1450_ = \o:n9->n10  & ~new_n1378_;
  assign new_n1451_ = ~\o:~n9->n10  & ~new_n1450_;
  assign new_n1452_ = ~\o:~n9->n70  & ~\o:n9->n71 ;
  assign new_n1453_ = ~\o:n9->n70  & new_n1452_;
  assign new_n1454_ = ~\o:~n9->n66  & new_n1453_;
  assign new_n1455_ = new_n1278_ & new_n1454_;
  assign new_n1456_ = ~\o:n9->n66  & new_n1455_;
  assign new_n1457_ = ~\o:~n9->n39  & new_n1456_;
  assign new_n1458_ = ~\o:n9->n39  & new_n1457_;
  assign new_n1459_ = ~\o:n9->n10  & new_n1374_;
  assign new_n1460_ = new_n1458_ & new_n1459_;
  assign new_n1461_ = ~new_n1451_ & ~new_n1460_;
  assign new_n1462_ = ~\o:~n9->n33  & new_n1154_;
  assign new_n1463_ = \o:n9->n33  & ~new_n1462_;
  assign new_n1464_ = ~\o:n68->n39  & new_n1044_;
  assign new_n1465_ = \o:~n68->n33  & ~new_n1464_;
  assign new_n1466_ = ~\o:n48->n4  & ~\o:~n48->n4 ;
  assign new_n1467_ = new_n992_ & new_n995_;
  assign new_n1468_ = \o:~n48->n4  & ~new_n1467_;
  assign new_n1469_ = new_n991_ & ~new_n1468_;
  assign new_n1470_ = ~new_n1466_ & ~new_n1469_;
  assign new_n1471_ = ~new_n1465_ & ~new_n1470_;
  assign new_n1472_ = ~new_n1463_ & new_n1471_;
  assign new_n1473_ = ~new_n1461_ & new_n1472_;
  assign new_n1474_ = \o:n65->n66  & ~new_n986_;
  assign new_n1475_ = \o:n56->n66  & ~new_n1032_;
  assign new_n1476_ = ~new_n1474_ & ~new_n1475_;
  assign new_n1477_ = ~\o:~n56->n66  & new_n1138_;
  assign new_n1478_ = ~\o:~n48->n66  & new_n1477_;
  assign new_n1479_ = ~\o:n56->n66  & new_n1478_;
  assign new_n1480_ = \o:n48->n66  & ~new_n1479_;
  assign new_n1481_ = new_n1160_ & new_n1205_;
  assign new_n1482_ = new_n1100_ & new_n1481_;
  assign new_n1483_ = ~new_n1161_ & ~new_n1482_;
  assign new_n1484_ = ~new_n1480_ & ~new_n1483_;
  assign new_n1485_ = \o:n65->n39  & ~new_n988_;
  assign new_n1486_ = ~\o:~n65->n4  & new_n1386_;
  assign new_n1487_ = \o:n65->n4  & ~new_n1486_;
  assign new_n1488_ = ~new_n1485_ & ~new_n1487_;
  assign new_n1489_ = ~\o:~n68->n4  & new_n1345_;
  assign new_n1490_ = \o:n68->n4  & ~new_n1489_;
  assign new_n1491_ = \o:n56->n39  & ~new_n1034_;
  assign new_n1492_ = ~new_n1490_ & ~new_n1491_;
  assign new_n1493_ = new_n1488_ & new_n1492_;
  assign new_n1494_ = new_n1484_ & new_n1493_;
  assign new_n1495_ = new_n1476_ & new_n1494_;
  assign new_n1496_ = new_n1473_ & new_n1495_;
  assign new_n1497_ = new_n1449_ & new_n1496_;
  assign new_n1498_ = ~\o:~n56->n4  & new_n992_;
  assign new_n1499_ = ~new_n991_ & ~new_n1498_;
  assign new_n1500_ = \o:n56->n71  & ~new_n1027_;
  assign new_n1501_ = ~\o:~n56->n70  & ~new_n1500_;
  assign new_n1502_ = ~new_n1060_ & ~new_n1501_;
  assign new_n1503_ = ~new_n1499_ & ~new_n1502_;
  assign new_n1504_ = \o:n77->n66  & ~new_n1182_;
  assign new_n1505_ = \o:n56->n10  & ~new_n1002_;
  assign new_n1506_ = new_n1001_ & ~new_n1505_;
  assign new_n1507_ = ~new_n1004_ & ~new_n1506_;
  assign new_n1508_ = ~\o:~n56->n4  & new_n993_;
  assign new_n1509_ = \o:n56->n4  & ~new_n1508_;
  assign new_n1510_ = ~new_n1507_ & ~new_n1509_;
  assign new_n1511_ = ~new_n1504_ & new_n1510_;
  assign new_n1512_ = new_n1503_ & new_n1511_;
  assign new_n1513_ = \o:~n9->n4  & ~new_n1380_;
  assign new_n1514_ = ~\o:n48->n70  & new_n1232_;
  assign new_n1515_ = ~\o:~n48->n66  & new_n1514_;
  assign new_n1516_ = new_n1227_ & new_n1515_;
  assign new_n1517_ = ~\o:n48->n66  & new_n1516_;
  assign new_n1518_ = ~\o:~n48->n39  & new_n1517_;
  assign new_n1519_ = ~\o:n48->n39  & new_n1518_;
  assign new_n1520_ = \o:~n48->n33  & ~new_n1519_;
  assign new_n1521_ = ~new_n1513_ & ~new_n1520_;
  assign new_n1522_ = new_n1512_ & new_n1521_;
  assign new_n1523_ = \o:n48->n39  & ~new_n1518_;
  assign new_n1524_ = \o:~n9->n33  & ~new_n1458_;
  assign new_n1525_ = ~new_n1523_ & ~new_n1524_;
  assign new_n1526_ = \o:~n48->n66  & ~new_n1443_;
  assign new_n1527_ = \o:n42->n39  & ~new_n1243_;
  assign new_n1528_ = ~\o:n48->n66  & ~\o:~n48->n71 ;
  assign new_n1529_ = new_n1515_ & new_n1528_;
  assign new_n1530_ = \o:~n48->n39  & ~new_n1529_;
  assign new_n1531_ = ~new_n1527_ & ~new_n1530_;
  assign new_n1532_ = ~new_n1526_ & new_n1531_;
  assign new_n1533_ = new_n1278_ & new_n1452_;
  assign new_n1534_ = ~\o:n9->n70  & new_n1533_;
  assign new_n1535_ = \o:~n9->n66  & ~new_n1534_;
  assign new_n1536_ = \o:n9->n70  & ~new_n1533_;
  assign new_n1537_ = \o:~n42->n39  & ~new_n1242_;
  assign new_n1538_ = ~new_n1536_ & ~new_n1537_;
  assign new_n1539_ = ~\o:n9->n66  & ~\o:~n9->n71 ;
  assign new_n1540_ = new_n1454_ & new_n1539_;
  assign new_n1541_ = \o:~n9->n39  & ~new_n1540_;
  assign new_n1542_ = new_n1538_ & ~new_n1541_;
  assign new_n1543_ = ~new_n1535_ & new_n1542_;
  assign new_n1544_ = new_n995_ & new_n1235_;
  assign new_n1545_ = new_n1061_ & new_n1544_;
  assign new_n1546_ = new_n992_ & new_n1389_;
  assign new_n1547_ = new_n1386_ & new_n1546_;
  assign new_n1548_ = ~new_n1545_ & ~new_n1547_;
  assign new_n1549_ = ~\o:~n68->n39  & new_n1204_;
  assign new_n1550_ = ~new_n1037_ & ~new_n1549_;
  assign new_n1551_ = ~\o:~n65->n39  & new_n1397_;
  assign new_n1552_ = ~new_n981_ & ~new_n1551_;
  assign new_n1553_ = ~new_n1550_ & ~new_n1552_;
  assign new_n1554_ = ~\o:~n42->n66  & ~\o:n42->n71 ;
  assign new_n1555_ = \o:~n42->n71  & ~new_n1554_;
  assign new_n1556_ = ~new_n1239_ & ~new_n1240_;
  assign new_n1557_ = \o:~n56->n39  & ~new_n1027_;
  assign new_n1558_ = ~new_n1556_ & ~new_n1557_;
  assign new_n1559_ = ~new_n1555_ & new_n1558_;
  assign new_n1560_ = new_n1553_ & new_n1559_;
  assign new_n1561_ = new_n1548_ & new_n1560_;
  assign new_n1562_ = new_n1543_ & new_n1561_;
  assign new_n1563_ = new_n1532_ & new_n1562_;
  assign new_n1564_ = new_n1525_ & new_n1563_;
  assign new_n1565_ = new_n1522_ & new_n1564_;
  assign new_n1566_ = new_n1497_ & new_n1565_;
  assign new_n1567_ = new_n1437_ & new_n1566_;
  assign new_n1568_ = ~\o:n48->n66  & new_n1479_;
  assign new_n1569_ = \o:~n42->n66  & ~new_n1568_;
  assign new_n1570_ = \o:n56->n66  & ~new_n1477_;
  assign new_n1571_ = ~\o:~n6->n70  & new_n1421_;
  assign new_n1572_ = \o:n6->n70  & ~new_n1571_;
  assign new_n1573_ = ~new_n1570_ & ~new_n1572_;
  assign new_n1574_ = new_n1072_ & new_n1077_;
  assign new_n1575_ = ~new_n1069_ & ~new_n1574_;
  assign new_n1576_ = ~\o:~n6->n66  & new_n1120_;
  assign new_n1577_ = \o:n6->n66  & ~new_n1576_;
  assign new_n1578_ = ~new_n1575_ & ~new_n1577_;
  assign new_n1579_ = new_n1573_ & new_n1578_;
  assign new_n1580_ = ~new_n1569_ & new_n1579_;
  assign new_n1581_ = \o:n48->n70  & ~new_n1024_;
  assign new_n1582_ = ~\o:~n9->n79  & new_n1113_;
  assign new_n1583_ = \o:n9->n79  & ~new_n1582_;
  assign new_n1584_ = \o:n56->n70  & ~new_n1022_;
  assign new_n1585_ = ~new_n1583_ & ~new_n1584_;
  assign new_n1586_ = ~new_n1581_ & new_n1585_;
  assign new_n1587_ = new_n1580_ & new_n1586_;
  assign new_n1588_ = new_n1118_ & new_n1568_;
  assign new_n1589_ = \o:~n9->n66  & ~new_n1588_;
  assign new_n1590_ = ~\o:n9->n66  & ~new_n1589_;
  assign new_n1591_ = ~\o:~n9->n66  & new_n1132_;
  assign new_n1592_ = new_n1120_ & new_n1591_;
  assign new_n1593_ = ~new_n1590_ & ~new_n1592_;
  assign new_n1594_ = new_n1151_ & new_n1464_;
  assign new_n1595_ = \o:~n68->n10  & ~new_n1594_;
  assign new_n1596_ = ~\o:n68->n10  & ~new_n1595_;
  assign new_n1597_ = ~\o:~n68->n10  & new_n1197_;
  assign new_n1598_ = new_n1345_ & new_n1597_;
  assign new_n1599_ = ~new_n1596_ & ~new_n1598_;
  assign new_n1600_ = new_n1000_ & new_n1445_;
  assign new_n1601_ = ~new_n1466_ & ~new_n1600_;
  assign new_n1602_ = new_n1441_ & new_n1519_;
  assign new_n1603_ = \o:~n48->n10  & ~new_n1602_;
  assign new_n1604_ = ~new_n1601_ & ~new_n1603_;
  assign new_n1605_ = ~new_n1599_ & new_n1604_;
  assign new_n1606_ = ~new_n1593_ & new_n1605_;
  assign new_n1607_ = new_n1587_ & new_n1606_;
  assign new_n1608_ = ~\o:n9->n70  & new_n1239_;
  assign new_n1609_ = new_n1025_ & new_n1608_;
  assign new_n1610_ = \o:~n9->n70  & ~new_n1609_;
  assign new_n1611_ = new_n989_ & new_n1144_;
  assign new_n1612_ = \o:~n65->n10  & ~new_n1611_;
  assign new_n1613_ = ~\o:n65->n10  & ~new_n1612_;
  assign new_n1614_ = ~\o:~n65->n10  & new_n1388_;
  assign new_n1615_ = new_n1386_ & new_n1614_;
  assign new_n1616_ = ~new_n1613_ & ~new_n1615_;
  assign new_n1617_ = ~new_n1610_ & ~new_n1616_;
  assign new_n1618_ = \o:n68->n70  & ~new_n1018_;
  assign new_n1619_ = ~\o:~n65->n70  & ~new_n1618_;
  assign new_n1620_ = ~new_n1415_ & ~new_n1619_;
  assign new_n1621_ = ~new_n1204_ & ~new_n1397_;
  assign new_n1622_ = new_n1097_ & ~new_n1621_;
  assign new_n1623_ = new_n1204_ & new_n1398_;
  assign new_n1624_ = ~new_n1622_ & ~new_n1623_;
  assign new_n1625_ = ~\o:~n56->n79  & new_n1037_;
  assign new_n1626_ = ~\o:~n56->n79  & new_n1226_;
  assign new_n1627_ = ~new_n1037_ & ~new_n1626_;
  assign new_n1628_ = new_n981_ & ~new_n1627_;
  assign new_n1629_ = ~new_n1625_ & ~new_n1628_;
  assign new_n1630_ = ~new_n1624_ & ~new_n1629_;
  assign new_n1631_ = ~new_n1620_ & new_n1630_;
  assign new_n1632_ = \o:n56->n79  & ~new_n1111_;
  assign new_n1633_ = \o:~n56->n4  & ~new_n992_;
  assign new_n1634_ = ~new_n1130_ & ~new_n1131_;
  assign new_n1635_ = ~\o:~n65->n66  & ~\o:~n68->n66 ;
  assign new_n1636_ = \o:n68->n66  & ~new_n1635_;
  assign new_n1637_ = ~new_n1634_ & ~new_n1636_;
  assign new_n1638_ = ~new_n1633_ & new_n1637_;
  assign new_n1639_ = ~\o:~n56->n33  & new_n1441_;
  assign new_n1640_ = ~new_n1151_ & ~new_n1639_;
  assign new_n1641_ = \o:n56->n33  & ~new_n1152_;
  assign new_n1642_ = ~new_n1640_ & ~new_n1641_;
  assign new_n1643_ = \o:~n65->n66  & ~new_n1135_;
  assign new_n1644_ = ~\o:~n56->n33  & new_n1151_;
  assign new_n1645_ = ~new_n1144_ & ~new_n1644_;
  assign new_n1646_ = ~new_n1643_ & ~new_n1645_;
  assign new_n1647_ = ~\o:n68->n70  & new_n1018_;
  assign new_n1648_ = \o:~n68->n70  & ~new_n1647_;
  assign new_n1649_ = ~\o:n56->n10  & new_n1002_;
  assign new_n1650_ = \o:~n56->n10  & ~new_n1649_;
  assign new_n1651_ = ~new_n1648_ & ~new_n1650_;
  assign new_n1652_ = new_n1646_ & new_n1651_;
  assign new_n1653_ = new_n1642_ & new_n1652_;
  assign new_n1654_ = new_n1638_ & new_n1653_;
  assign new_n1655_ = ~new_n1632_ & new_n1654_;
  assign new_n1656_ = new_n1631_ & new_n1655_;
  assign new_n1657_ = \o:n9->n4  & ~new_n1381_;
  assign new_n1658_ = \o:n48->n66  & ~new_n1516_;
  assign new_n1659_ = \o:n9->n39  & ~new_n1457_;
  assign new_n1660_ = ~new_n1658_ & ~new_n1659_;
  assign new_n1661_ = ~new_n1657_ & new_n1660_;
  assign new_n1662_ = ~\o:~n56->n4  & new_n1061_;
  assign new_n1663_ = \o:n56->n4  & ~new_n1662_;
  assign new_n1664_ = \o:n9->n66  & ~new_n1455_;
  assign new_n1665_ = ~new_n1663_ & ~new_n1664_;
  assign new_n1666_ = new_n1466_ & new_n1600_;
  assign new_n1667_ = ~\o:~n9->n33  & new_n1533_;
  assign new_n1668_ = ~\o:n9->n70  & new_n1375_;
  assign new_n1669_ = new_n1129_ & new_n1668_;
  assign new_n1670_ = new_n1667_ & new_n1669_;
  assign new_n1671_ = \o:n9->n33  & ~new_n1670_;
  assign new_n1672_ = ~new_n1666_ & ~new_n1671_;
  assign new_n1673_ = new_n991_ & new_n1345_;
  assign new_n1674_ = new_n1198_ & new_n1673_;
  assign new_n1675_ = \o:~n48->n70  & ~new_n1018_;
  assign new_n1676_ = ~\o:~n65->n39  & ~\o:~n77->n39 ;
  assign new_n1677_ = \o:n65->n39  & ~new_n1676_;
  assign new_n1678_ = ~new_n1071_ & ~new_n1088_;
  assign new_n1679_ = \o:~n48->n66  & ~new_n1131_;
  assign new_n1680_ = ~new_n1678_ & ~new_n1679_;
  assign new_n1681_ = ~new_n1677_ & new_n1680_;
  assign new_n1682_ = ~new_n1675_ & new_n1681_;
  assign new_n1683_ = ~\o:~n48->n39  & new_n1160_;
  assign new_n1684_ = ~new_n1226_ & ~new_n1683_;
  assign new_n1685_ = new_n1128_ & new_n1328_;
  assign new_n1686_ = \o:~n9->n39  & ~new_n1277_;
  assign new_n1687_ = ~new_n1685_ & ~new_n1686_;
  assign new_n1688_ = ~\o:n42->n4  & ~\o:~n42->n79 ;
  assign new_n1689_ = ~\o:n42->n79  & new_n1688_;
  assign new_n1690_ = ~\o:n42->n10  & ~\o:~n42->n10 ;
  assign new_n1691_ = ~\o:~n42->n4  & new_n1690_;
  assign new_n1692_ = new_n1689_ & new_n1691_;
  assign new_n1693_ = new_n1687_ & new_n1692_;
  assign new_n1694_ = ~new_n1684_ & new_n1693_;
  assign new_n1695_ = ~\o:n42->n33  & ~\o:~n42->n33 ;
  assign new_n1696_ = ~\o:n77->n10  & ~\o:~n77->n10 ;
  assign new_n1697_ = new_n1695_ & new_n1696_;
  assign new_n1698_ = ~\o:n65->n39  & ~\o:~n77->n39 ;
  assign new_n1699_ = \o:n77->n39  & ~new_n1698_;
  assign new_n1700_ = ~\o:n77->n33  & ~\o:~n77->n33 ;
  assign new_n1701_ = ~\o:n77->n79  & ~\o:~n77->n79 ;
  assign new_n1702_ = ~\o:n77->n4  & ~\o:~n77->n4 ;
  assign new_n1703_ = new_n1701_ & new_n1702_;
  assign new_n1704_ = new_n1700_ & new_n1703_;
  assign new_n1705_ = ~new_n1699_ & new_n1704_;
  assign new_n1706_ = new_n1697_ & new_n1705_;
  assign new_n1707_ = new_n1694_ & new_n1706_;
  assign new_n1708_ = new_n1682_ & new_n1707_;
  assign new_n1709_ = ~new_n1674_ & new_n1708_;
  assign new_n1710_ = new_n1672_ & new_n1709_;
  assign new_n1711_ = new_n1665_ & new_n1710_;
  assign new_n1712_ = new_n1661_ & new_n1711_;
  assign new_n1713_ = new_n1656_ & new_n1712_;
  assign new_n1714_ = new_n1617_ & new_n1713_;
  assign new_n1715_ = new_n1607_ & new_n1714_;
  assign new_n1716_ = new_n1567_ & new_n1715_;
  assign new_n1717_ = ~new_n980_ & new_n1716_;
  assign new_n1718_ = ~new_n979_ & new_n1717_;
  assign new_n1719_ = new_n975_ & new_n1718_;
  assign new_n1720_ = new_n969_ & new_n1719_;
  assign new_n1721_ = ~new_n966_ & new_n1720_;
  assign new_n1722_ = new_n960_ & new_n1721_;
  assign new_n1723_ = new_n716_ & ~new_n756_;
  assign new_n1724_ = ~new_n716_ & new_n756_;
  assign new_n1725_ = ~new_n1723_ & ~new_n1724_;
  assign new_n1726_ = \o:~n6->n70  & new_n1725_;
  assign new_n1727_ = \o:n6->n70  & ~new_n1725_;
  assign new_n1728_ = ~new_n1726_ & ~new_n1727_;
  assign new_n1729_ = \o:~n42->n71  & new_n856_;
  assign new_n1730_ = new_n708_ & ~new_n756_;
  assign new_n1731_ = ~new_n708_ & new_n756_;
  assign new_n1732_ = ~new_n1730_ & ~new_n1731_;
  assign new_n1733_ = \o:~n6->n66  & new_n1732_;
  assign new_n1734_ = \o:n6->n66  & ~new_n1732_;
  assign new_n1735_ = ~new_n1733_ & ~new_n1734_;
  assign new_n1736_ = ~new_n1729_ & new_n1735_;
  assign new_n1737_ = new_n1728_ & new_n1736_;
  assign new_n1738_ = ~new_n715_ & ~new_n751_;
  assign new_n1739_ = new_n715_ & new_n751_;
  assign new_n1740_ = ~new_n1738_ & ~new_n1739_;
  assign new_n1741_ = ~\o:~n9->n4  & new_n1740_;
  assign new_n1742_ = ~\o:n9->n4  & ~new_n1740_;
  assign new_n1743_ = ~new_n1741_ & ~new_n1742_;
  assign new_n1744_ = new_n1737_ & ~new_n1743_;
  assign new_n1745_ = ~new_n686_ & ~new_n715_;
  assign new_n1746_ = new_n686_ & new_n715_;
  assign new_n1747_ = ~new_n1745_ & ~new_n1746_;
  assign new_n1748_ = \o:n68->n4  & ~new_n1747_;
  assign new_n1749_ = \o:~n68->n4  & new_n1747_;
  assign new_n1750_ = ~new_n1748_ & ~new_n1749_;
  assign new_n1751_ = ~new_n708_ & ~new_n751_;
  assign new_n1752_ = new_n708_ & new_n751_;
  assign new_n1753_ = ~new_n1751_ & ~new_n1752_;
  assign new_n1754_ = ~\o:~n9->n66  & new_n1753_;
  assign new_n1755_ = ~\o:n9->n66  & ~new_n1753_;
  assign new_n1756_ = ~new_n1754_ & ~new_n1755_;
  assign new_n1757_ = new_n1750_ & ~new_n1756_;
  assign new_n1758_ = new_n1744_ & new_n1757_;
  assign new_n1759_ = new_n1722_ & new_n1758_;
  assign new_n1760_ = ~new_n947_ & new_n1759_;
  assign new_n1761_ = ~new_n246_ & new_n772_;
  assign new_n1762_ = new_n246_ & ~new_n772_;
  assign new_n1763_ = ~new_n1761_ & ~new_n1762_;
  assign new_n1764_ = \o:n56->n33  & ~new_n1763_;
  assign new_n1765_ = \o:~n56->n33  & new_n1763_;
  assign new_n1766_ = ~new_n1764_ & ~new_n1765_;
  assign new_n1767_ = new_n1760_ & new_n1766_;
  assign new_n1768_ = new_n943_ & new_n1767_;
  assign new_n1769_ = new_n930_ & new_n1768_;
  assign new_n1770_ = new_n870_ & new_n1769_;
  assign new_n1771_ = new_n246_ & ~new_n787_;
  assign new_n1772_ = ~new_n1761_ & ~new_n1771_;
  assign new_n1773_ = \o:n56->n10  & new_n1772_;
  assign new_n1774_ = \o:~n56->n10  & ~new_n1772_;
  assign new_n1775_ = ~new_n652_ & ~new_n693_;
  assign new_n1776_ = new_n652_ & new_n693_;
  assign new_n1777_ = ~new_n1775_ & ~new_n1776_;
  assign new_n1778_ = new_n246_ & ~new_n1777_;
  assign new_n1779_ = ~new_n876_ & ~new_n1778_;
  assign new_n1780_ = \o:n48->n10  & new_n1779_;
  assign new_n1781_ = \o:~n48->n10  & ~new_n1779_;
  assign new_n1782_ = new_n652_ & ~new_n718_;
  assign new_n1783_ = ~new_n652_ & new_n718_;
  assign new_n1784_ = ~new_n1782_ & ~new_n1783_;
  assign new_n1785_ = \o:n48->n79  & ~new_n1784_;
  assign new_n1786_ = \o:~n48->n79  & new_n1784_;
  assign new_n1787_ = ~new_n1785_ & ~new_n1786_;
  assign new_n1788_ = ~\o:~n48->n71  & new_n1777_;
  assign new_n1789_ = ~\o:n48->n71  & ~new_n1777_;
  assign new_n1790_ = ~new_n1788_ & ~new_n1789_;
  assign new_n1791_ = new_n1787_ & ~new_n1790_;
  assign new_n1792_ = ~new_n1781_ & new_n1791_;
  assign new_n1793_ = ~new_n1780_ & new_n1792_;
  assign new_n1794_ = ~new_n1774_ & new_n1793_;
  assign new_n1795_ = ~new_n1773_ & new_n1794_;
  assign new_n1796_ = new_n652_ & ~new_n715_;
  assign new_n1797_ = ~new_n652_ & new_n715_;
  assign new_n1798_ = ~new_n1796_ & ~new_n1797_;
  assign new_n1799_ = \o:n48->n4  & ~new_n1798_;
  assign new_n1800_ = \o:~n48->n4  & new_n1798_;
  assign new_n1801_ = ~new_n1799_ & ~new_n1800_;
  assign new_n1802_ = ~new_n686_ & ~new_n716_;
  assign new_n1803_ = new_n686_ & new_n716_;
  assign new_n1804_ = ~new_n1802_ & ~new_n1803_;
  assign new_n1805_ = ~\o:~n68->n70  & new_n1804_;
  assign new_n1806_ = ~\o:n68->n70  & ~new_n1804_;
  assign new_n1807_ = ~new_n1805_ & ~new_n1806_;
  assign new_n1808_ = ~\o:~n68->n71  & new_n696_;
  assign new_n1809_ = ~\o:n68->n71  & ~new_n696_;
  assign new_n1810_ = ~new_n1808_ & ~new_n1809_;
  assign new_n1811_ = ~new_n1807_ & ~new_n1810_;
  assign new_n1812_ = new_n1801_ & new_n1811_;
  assign new_n1813_ = ~new_n715_ & ~new_n764_;
  assign new_n1814_ = new_n715_ & new_n764_;
  assign new_n1815_ = ~new_n1813_ & ~new_n1814_;
  assign new_n1816_ = \o:n65->n4  & ~new_n1815_;
  assign new_n1817_ = new_n246_ & new_n956_;
  assign new_n1818_ = ~new_n884_ & ~new_n1817_;
  assign new_n1819_ = \o:~n9->n10  & new_n1818_;
  assign new_n1820_ = ~new_n1816_ & ~new_n1819_;
  assign new_n1821_ = \o:n9->n10  & ~new_n1818_;
  assign new_n1822_ = ~new_n704_ & ~new_n764_;
  assign new_n1823_ = new_n704_ & new_n764_;
  assign new_n1824_ = ~new_n1822_ & ~new_n1823_;
  assign new_n1825_ = \o:n65->n39  & ~new_n1824_;
  assign new_n1826_ = \o:~n65->n39  & new_n1824_;
  assign new_n1827_ = ~new_n1825_ & ~new_n1826_;
  assign new_n1828_ = ~new_n1821_ & new_n1827_;
  assign new_n1829_ = new_n1820_ & new_n1828_;
  assign new_n1830_ = new_n1812_ & new_n1829_;
  assign new_n1831_ = \o:n56->n70  & ~new_n783_;
  assign new_n1832_ = \o:~n56->n4  & new_n946_;
  assign new_n1833_ = ~new_n1831_ & ~new_n1832_;
  assign new_n1834_ = \o:~n65->n4  & new_n1815_;
  assign new_n1835_ = \o:n65->n33  & new_n925_;
  assign new_n1836_ = ~new_n1834_ & ~new_n1835_;
  assign new_n1837_ = new_n246_ & new_n917_;
  assign new_n1838_ = ~new_n923_ & ~new_n1837_;
  assign new_n1839_ = \o:~n65->n10  & new_n1838_;
  assign new_n1840_ = \o:n65->n10  & ~new_n1838_;
  assign new_n1841_ = ~new_n1839_ & ~new_n1840_;
  assign new_n1842_ = new_n1836_ & new_n1841_;
  assign new_n1843_ = new_n1833_ & new_n1842_;
  assign new_n1844_ = new_n1830_ & new_n1843_;
  assign new_n1845_ = new_n1795_ & new_n1844_;
  assign n4381 = new_n1770_ & new_n1845_;
endmodule


